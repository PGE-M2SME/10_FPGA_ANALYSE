// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.3.469
// Netlist written on Mon Mar 29 18:33:38 2021
//
// Verilog Description of module test_DVI
//

module test_DVI (DE, Vsync, Hsync, ODCK, Hdisp, Vdisp, Hblank, 
            Vblank, Hsync_out, Vsync_out);   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(36[8:16])
    input DE;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(39[1:3])
    input Vsync;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(40[1:6])
    input Hsync;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(41[1:6])
    input ODCK;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(42[1:5])
    output [15:0]Hdisp;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    output [15:0]Vdisp;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    output [15:0]Hblank;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    output [15:0]Vblank;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    output [15:0]Hsync_out;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    output [15:0]Vsync_out;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    
    wire ODCK_c /* synthesis SET_AS_NETWORK=ODCK_c, is_clock=1 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(42[1:5])
    
    wire GND_net, VCC_net, DE_c, Vsync_c, Hsync_c, Hdisp_c_15, Hdisp_c_14, 
        Hdisp_c_13, Hdisp_c_12, Hdisp_c_11, Hdisp_c_10, Hdisp_c_9, 
        Hdisp_c_8, Hdisp_c_7, Hdisp_c_6, Hdisp_c_5, Hdisp_c_4, Hdisp_c_3, 
        Hdisp_c_2, Hdisp_c_1, Hdisp_c_0, Vdisp_c_15, Vdisp_c_14, Vdisp_c_13, 
        Vdisp_c_12, Vdisp_c_11, Vdisp_c_10, Vdisp_c_9, Vdisp_c_8, 
        Vdisp_c_7, Vdisp_c_6, Vdisp_c_5, Vdisp_c_4, Vdisp_c_3, Vdisp_c_2, 
        Vdisp_c_1, Vdisp_c_0, Hblank_c_15, Hblank_c_14, Hblank_c_13, 
        Hblank_c_12, Hblank_c_11, Hblank_c_10, Hblank_c_9, Hblank_c_8, 
        Hblank_c_7, Hblank_c_6, Hblank_c_5, Hblank_c_4, Hblank_c_3, 
        Hblank_c_2, Hblank_c_1, Hblank_c_0, Vblank_c_15, Vblank_c_14, 
        Vblank_c_13, Vblank_c_12, Vblank_c_11, Vblank_c_10, Vblank_c_9, 
        Vblank_c_8, Vblank_c_7, Vblank_c_6, Vblank_c_5, Vblank_c_4, 
        Vblank_c_3, Vblank_c_2, Vblank_c_1, Vblank_c_0, Hsync_out_c_15, 
        Hsync_out_c_14, Hsync_out_c_13, Hsync_out_c_12, Hsync_out_c_11, 
        Hsync_out_c_10, Hsync_out_c_9, Hsync_out_c_8, Hsync_out_c_7, 
        Hsync_out_c_6, Hsync_out_c_5, Hsync_out_c_4, Hsync_out_c_3, 
        Hsync_out_c_2, Hsync_out_c_1, Hsync_out_c_0, Vsync_out_c_15, 
        Vsync_out_c_14, Vsync_out_c_13, Vsync_out_c_12, Vsync_out_c_11, 
        Vsync_out_c_10, Vsync_out_c_9, Vsync_out_c_8, Vsync_out_c_7, 
        Vsync_out_c_6, Vsync_out_c_5, Vsync_out_c_4, Vsync_out_c_3, 
        Vsync_out_c_2, Vsync_out_c_1, Vsync_out_c_0;
    wire [15:0]sig_Hdisp_cpt;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(56[8:21])
    wire [15:0]sig_compt_front_Hsync;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(63[8:29])
    
    wire out_comp, rising_Hsync, detect, D_detect, detect_DE, D_detect_DE, 
        n1263, ODCK_c_enable_96, n1262, n1296, n1295, n1294, n1257, 
        n1259, n85, n84, n83, n82, n81, n80, n79, n78, n77, 
        n76, n75, n74, n73, n26, n22, n85_adj_1, n84_adj_2, 
        n83_adj_3, n82_adj_4, n81_adj_5, n80_adj_6, n79_adj_7, n78_adj_8, 
        n77_adj_9, n76_adj_10, n75_adj_11, n74_adj_12, n73_adj_13, 
        n72, n71, n70, n1261, n72_adj_14, n71_adj_15, n70_adj_16, 
        n20, n30, n28, n18, n17, n1281, n85_adj_17, n84_adj_18, 
        n31, n29, n83_adj_19, n82_adj_20, n81_adj_21, n80_adj_22, 
        n79_adj_23, n78_adj_24, n77_adj_25, n76_adj_26, n75_adj_27, 
        n74_adj_28, n73_adj_29, n72_adj_30, n71_adj_31, n70_adj_32, 
        n1256, n1264, n1260, out_comp_N_378, n1292, n1291, n1290, 
        n1289, n1288, n1285, n1284, n1282, n1084, n1258, n1297, 
        n70_adj_33, n71_adj_34, n72_adj_35, n73_adj_36, n74_adj_37, 
        n75_adj_38, n76_adj_39, n77_adj_40, n78_adj_41, n79_adj_42, 
        n80_adj_43, n81_adj_44, n82_adj_45, n83_adj_46, n84_adj_47, 
        n85_adj_48, n70_adj_49, n71_adj_50, n72_adj_51, n73_adj_52, 
        n74_adj_53, n75_adj_54, n76_adj_55, n77_adj_56, n78_adj_57, 
        n79_adj_58, n80_adj_59, n81_adj_60, n82_adj_61, n83_adj_62, 
        n84_adj_63, n85_adj_64, n28_adj_65, n1114, ODCK_c_enable_92, 
        n26_adj_66, n25, n1381, ODCK_c_enable_97, n1293, n1283, 
        ODCK_c_enable_95, n70_adj_67, n71_adj_68, n72_adj_69, n73_adj_70, 
        n74_adj_71, n75_adj_72, n76_adj_73, n77_adj_74, n78_adj_75, 
        n79_adj_76, n80_adj_77, n81_adj_78, n82_adj_79, n83_adj_80, 
        n84_adj_81, n85_adj_82, n1280, n1298, n1278, n1277, n1276, 
        n1275, n1274, n1273, n1272, n1271, n1270, n1269, n1268, 
        n1267, n1266, n1310, ODCK_c_enable_94, n1286, ODCK_c_enable_93, 
        n70_adj_83, n71_adj_84, n72_adj_85, n73_adj_86, n74_adj_87, 
        n75_adj_88, n76_adj_89, n77_adj_90, n78_adj_91, n79_adj_92, 
        n80_adj_93, n81_adj_94, n82_adj_95, n83_adj_96, n84_adj_97, 
        n85_adj_98, n1309, n1308, n1307, n1306, n1305, n1304, 
        n1303, n1302, n1301, n1300, n1299, n1265, n1279, n1311, 
        n1380, ODCK_c_enable_17, n1287;
    
    VHI i2 (.Z(VCC_net));
    OB Hdisp_pad_8 (.I(Hdisp_c_8), .O(Hdisp[8]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    CCU2C sig_compt_front_Hsync_156_add_4_17 (.A0(sig_compt_front_Hsync[15]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n1263), .S0(n70_adj_32));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156_add_4_17.INIT0 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_17.INIT1 = 16'h0000;
    defparam sig_compt_front_Hsync_156_add_4_17.INJECT1_0 = "NO";
    defparam sig_compt_front_Hsync_156_add_4_17.INJECT1_1 = "NO";
    OB Hdisp_pad_9 (.I(Hdisp_c_9), .O(Hdisp[9]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    FD1P3IX sig_compt_front_Hsync_156__i0 (.D(n85_adj_17), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i0.GSR = "ENABLED";
    CCU2C sig_compt_front_Hsync_156_add_4_1 (.A0(GND_net), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(sig_compt_front_Hsync[0]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .COUT(n1256), .S1(n85_adj_17));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156_add_4_1.INIT0 = 16'h0000;
    defparam sig_compt_front_Hsync_156_add_4_1.INIT1 = 16'h555f;
    defparam sig_compt_front_Hsync_156_add_4_1.INJECT1_0 = "NO";
    defparam sig_compt_front_Hsync_156_add_4_1.INJECT1_1 = "NO";
    CCU2C sig_compt_front_Hsync_156_add_4_3 (.A0(sig_compt_front_Hsync[1]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(sig_compt_front_Hsync[2]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n1256), .COUT(n1257), 
          .S0(n84_adj_18), .S1(n83_adj_19));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156_add_4_3.INIT0 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_3.INIT1 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_3.INJECT1_0 = "NO";
    defparam sig_compt_front_Hsync_156_add_4_3.INJECT1_1 = "NO";
    CCU2C sig_compt_front_Hsync_156_add_4_7 (.A0(sig_compt_front_Hsync[5]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(sig_compt_front_Hsync[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n1258), .COUT(n1259), 
          .S0(n80_adj_22), .S1(n79_adj_23));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156_add_4_7.INIT0 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_7.INIT1 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_7.INJECT1_0 = "NO";
    defparam sig_compt_front_Hsync_156_add_4_7.INJECT1_1 = "NO";
    CCU2C sig_compt_front_Hsync_156_add_4_15 (.A0(sig_compt_front_Hsync[13]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(sig_compt_front_Hsync[14]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n1262), .COUT(n1263), 
          .S0(n72_adj_30), .S1(n71_adj_31));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156_add_4_15.INIT0 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_15.INIT1 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_15.INJECT1_0 = "NO";
    defparam sig_compt_front_Hsync_156_add_4_15.INJECT1_1 = "NO";
    OB Hdisp_pad_10 (.I(Hdisp_c_10), .O(Hdisp[10]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    LUT4 i8_2_lut (.A(sig_compt_front_Hsync[2]), .B(sig_compt_front_Hsync[7]), 
         .Z(n25)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut.init = 16'heeee;
    FD1P3AX sig_Hdisp_i0_i1 (.D(sig_Hdisp_cpt[0]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_0)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i1.GSR = "ENABLED";
    CCU2C sig_Hsync_151_add_4_17 (.A0(Hsync_out_c_15), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n1295), .S0(n70_adj_49));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151_add_4_17.INIT0 = 16'haaa0;
    defparam sig_Hsync_151_add_4_17.INIT1 = 16'h0000;
    defparam sig_Hsync_151_add_4_17.INJECT1_0 = "NO";
    defparam sig_Hsync_151_add_4_17.INJECT1_1 = "NO";
    FD1S3AX detect_91 (.D(Hsync_c), .CK(ODCK_c), .Q(detect)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(183[1] 186[10])
    defparam detect_91.GSR = "ENABLED";
    OB Hdisp_pad_11 (.I(Hdisp_c_11), .O(Hdisp[11]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    GSR GSR_INST (.GSR(VCC_net));
    OB Hdisp_pad_12 (.I(Hdisp_c_12), .O(Hdisp[12]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    FD1S3AX D_detect_92 (.D(detect), .CK(ODCK_c), .Q(D_detect)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(183[1] 186[10])
    defparam D_detect_92.GSR = "ENABLED";
    FD1S3AX detect_DE_93 (.D(DE_c), .CK(ODCK_c), .Q(detect_DE)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(196[1] 199[10])
    defparam detect_DE_93.GSR = "ENABLED";
    FD1S3AX D_detect_DE_94 (.D(detect_DE), .CK(ODCK_c), .Q(D_detect_DE)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(196[1] 199[10])
    defparam D_detect_DE_94.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i1 (.D(n85), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_0)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i1.GSR = "ENABLED";
    CCU2C sig_Hblank_154_add_4_15 (.A0(Hblank_c_13), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hblank_c_14), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1278), .COUT(n1279), .S0(n72_adj_14), 
          .S1(n71_adj_15));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154_add_4_15.INIT0 = 16'haaa0;
    defparam sig_Hblank_154_add_4_15.INIT1 = 16'haaa0;
    defparam sig_Hblank_154_add_4_15.INJECT1_0 = "NO";
    defparam sig_Hblank_154_add_4_15.INJECT1_1 = "NO";
    OB Hdisp_pad_13 (.I(Hdisp_c_13), .O(Hdisp[13]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    CCU2C sig_compt_front_Hsync_156_add_4_13 (.A0(sig_compt_front_Hsync[11]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(sig_compt_front_Hsync[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n1261), .COUT(n1262), 
          .S0(n74_adj_28), .S1(n73_adj_29));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156_add_4_13.INIT0 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_13.INIT1 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_13.INJECT1_0 = "NO";
    defparam sig_compt_front_Hsync_156_add_4_13.INJECT1_1 = "NO";
    CCU2C sig_compt_front_Hsync_156_add_4_5 (.A0(sig_compt_front_Hsync[3]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(sig_compt_front_Hsync[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n1257), .COUT(n1258), 
          .S0(n82_adj_20), .S1(n81_adj_21));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156_add_4_5.INIT0 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_5.INIT1 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_5.INJECT1_0 = "NO";
    defparam sig_compt_front_Hsync_156_add_4_5.INJECT1_1 = "NO";
    CCU2C sig_Hblank_154_add_4_13 (.A0(Hblank_c_11), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hblank_c_12), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1277), .COUT(n1278), .S0(n74), .S1(n73));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154_add_4_13.INIT0 = 16'haaa0;
    defparam sig_Hblank_154_add_4_13.INIT1 = 16'haaa0;
    defparam sig_Hblank_154_add_4_13.INJECT1_0 = "NO";
    defparam sig_Hblank_154_add_4_13.INJECT1_1 = "NO";
    CCU2C sig_Hsync_151_add_4_15 (.A0(Hsync_out_c_13), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hsync_out_c_14), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1294), .COUT(n1295), .S0(n72_adj_51), 
          .S1(n71_adj_50));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151_add_4_15.INIT0 = 16'haaa0;
    defparam sig_Hsync_151_add_4_15.INIT1 = 16'haaa0;
    defparam sig_Hsync_151_add_4_15.INJECT1_0 = "NO";
    defparam sig_Hsync_151_add_4_15.INJECT1_1 = "NO";
    OB Hdisp_pad_14 (.I(Hdisp_c_14), .O(Hdisp[14]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    OB Hdisp_pad_15 (.I(Hdisp_c_15), .O(Hdisp[15]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    CCU2C sig_Hblank_154_add_4_11 (.A0(Hblank_c_9), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hblank_c_10), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1276), .COUT(n1277), .S0(n76), .S1(n75));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154_add_4_11.INIT0 = 16'haaa0;
    defparam sig_Hblank_154_add_4_11.INIT1 = 16'haaa0;
    defparam sig_Hblank_154_add_4_11.INJECT1_0 = "NO";
    defparam sig_Hblank_154_add_4_11.INJECT1_1 = "NO";
    CCU2C sig_Hblank_154_add_4_9 (.A0(Hblank_c_7), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hblank_c_8), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1275), .COUT(n1276), .S0(n78), .S1(n77));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154_add_4_9.INIT0 = 16'haaa0;
    defparam sig_Hblank_154_add_4_9.INIT1 = 16'haaa0;
    defparam sig_Hblank_154_add_4_9.INJECT1_0 = "NO";
    defparam sig_Hblank_154_add_4_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(DE_c), .B(Vsync_c), .C(detect_DE), .D(D_detect_DE), 
         .Z(ODCK_c_enable_93)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B+!(C+!(D))))) */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(39[1:3])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h4f44;
    CCU2C sig_Hdisp_cpt_147_add_4_7 (.A0(sig_Hdisp_cpt[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(sig_Hdisp_cpt[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n1306), .COUT(n1307), .S0(n80_adj_93), 
          .S1(n79_adj_92));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147_add_4_7.INIT0 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_7.INIT1 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_7.INJECT1_0 = "NO";
    defparam sig_Hdisp_cpt_147_add_4_7.INJECT1_1 = "NO";
    LUT4 i9_3_lut (.A(sig_compt_front_Hsync[1]), .B(DE_c), .C(sig_compt_front_Hsync[0]), 
         .Z(n26_adj_66)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i9_3_lut.init = 16'hfefe;
    LUT4 i70_2_lut_rep_6 (.A(out_comp), .B(DE_c), .Z(n1381)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(173[9:35])
    defparam i70_2_lut_rep_6.init = 16'h4444;
    CCU2C sig_Hblank_154_add_4_7 (.A0(Hblank_c_5), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hblank_c_6), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1274), .COUT(n1275), .S0(n80), .S1(n79));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154_add_4_7.INIT0 = 16'haaa0;
    defparam sig_Hblank_154_add_4_7.INIT1 = 16'haaa0;
    defparam sig_Hblank_154_add_4_7.INJECT1_0 = "NO";
    defparam sig_Hblank_154_add_4_7.INJECT1_1 = "NO";
    CCU2C sig_Hblank_154_add_4_5 (.A0(Hblank_c_3), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hblank_c_4), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1273), .COUT(n1274), .S0(n82), .S1(n81));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154_add_4_5.INIT0 = 16'haaa0;
    defparam sig_Hblank_154_add_4_5.INIT1 = 16'haaa0;
    defparam sig_Hblank_154_add_4_5.INJECT1_0 = "NO";
    defparam sig_Hblank_154_add_4_5.INJECT1_1 = "NO";
    CCU2C sig_Hblank_154_add_4_3 (.A0(Hblank_c_1), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hblank_c_2), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1272), .COUT(n1273), .S0(n84), .S1(n83));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154_add_4_3.INIT0 = 16'haaa0;
    defparam sig_Hblank_154_add_4_3.INIT1 = 16'haaa0;
    defparam sig_Hblank_154_add_4_3.INJECT1_0 = "NO";
    defparam sig_Hblank_154_add_4_3.INJECT1_1 = "NO";
    CCU2C sig_Hblank_154_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Hblank_c_0), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n1272), .S1(n85));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154_add_4_1.INIT0 = 16'h0000;
    defparam sig_Hblank_154_add_4_1.INIT1 = 16'h555f;
    defparam sig_Hblank_154_add_4_1.INJECT1_0 = "NO";
    defparam sig_Hblank_154_add_4_1.INJECT1_1 = "NO";
    CCU2C sig_Vblank_158_add_4_17 (.A0(Vblank_c_15), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n1271), .S0(n70));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158_add_4_17.INIT0 = 16'haaa0;
    defparam sig_Vblank_158_add_4_17.INIT1 = 16'h0000;
    defparam sig_Vblank_158_add_4_17.INJECT1_0 = "NO";
    defparam sig_Vblank_158_add_4_17.INJECT1_1 = "NO";
    CCU2C sig_Vblank_158_add_4_15 (.A0(Vblank_c_13), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vblank_c_14), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1270), .COUT(n1271), .S0(n72), .S1(n71));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158_add_4_15.INIT0 = 16'haaa0;
    defparam sig_Vblank_158_add_4_15.INIT1 = 16'haaa0;
    defparam sig_Vblank_158_add_4_15.INJECT1_0 = "NO";
    defparam sig_Vblank_158_add_4_15.INJECT1_1 = "NO";
    CCU2C sig_Vblank_158_add_4_13 (.A0(Vblank_c_11), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vblank_c_12), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1269), .COUT(n1270), .S0(n74_adj_12), 
          .S1(n73_adj_13));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158_add_4_13.INIT0 = 16'haaa0;
    defparam sig_Vblank_158_add_4_13.INIT1 = 16'haaa0;
    defparam sig_Vblank_158_add_4_13.INJECT1_0 = "NO";
    defparam sig_Vblank_158_add_4_13.INJECT1_1 = "NO";
    CCU2C sig_Vblank_158_add_4_11 (.A0(Vblank_c_9), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vblank_c_10), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1268), .COUT(n1269), .S0(n76_adj_10), 
          .S1(n75_adj_11));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158_add_4_11.INIT0 = 16'haaa0;
    defparam sig_Vblank_158_add_4_11.INIT1 = 16'haaa0;
    defparam sig_Vblank_158_add_4_11.INJECT1_0 = "NO";
    defparam sig_Vblank_158_add_4_11.INJECT1_1 = "NO";
    CCU2C sig_Vblank_158_add_4_9 (.A0(Vblank_c_7), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vblank_c_8), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1267), .COUT(n1268), .S0(n78_adj_8), .S1(n77_adj_9));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158_add_4_9.INIT0 = 16'haaa0;
    defparam sig_Vblank_158_add_4_9.INIT1 = 16'haaa0;
    defparam sig_Vblank_158_add_4_9.INJECT1_0 = "NO";
    defparam sig_Vblank_158_add_4_9.INJECT1_1 = "NO";
    CCU2C sig_Vblank_158_add_4_7 (.A0(Vblank_c_5), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vblank_c_6), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1266), .COUT(n1267), .S0(n80_adj_6), .S1(n79_adj_7));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158_add_4_7.INIT0 = 16'haaa0;
    defparam sig_Vblank_158_add_4_7.INIT1 = 16'haaa0;
    defparam sig_Vblank_158_add_4_7.INJECT1_0 = "NO";
    defparam sig_Vblank_158_add_4_7.INJECT1_1 = "NO";
    CCU2C sig_Vblank_158_add_4_5 (.A0(Vblank_c_3), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vblank_c_4), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1265), .COUT(n1266), .S0(n82_adj_4), .S1(n81_adj_5));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158_add_4_5.INIT0 = 16'haaa0;
    defparam sig_Vblank_158_add_4_5.INIT1 = 16'haaa0;
    defparam sig_Vblank_158_add_4_5.INJECT1_0 = "NO";
    defparam sig_Vblank_158_add_4_5.INJECT1_1 = "NO";
    CCU2C sig_Vblank_158_add_4_3 (.A0(Vblank_c_1), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vblank_c_2), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1264), .COUT(n1265), .S0(n84_adj_2), .S1(n83_adj_3));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158_add_4_3.INIT0 = 16'haaa0;
    defparam sig_Vblank_158_add_4_3.INIT1 = 16'haaa0;
    defparam sig_Vblank_158_add_4_3.INJECT1_0 = "NO";
    defparam sig_Vblank_158_add_4_3.INJECT1_1 = "NO";
    CCU2C sig_Vblank_158_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Vblank_c_0), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n1264), .S1(n85_adj_1));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158_add_4_1.INIT0 = 16'h0000;
    defparam sig_Vblank_158_add_4_1.INIT1 = 16'h555f;
    defparam sig_Vblank_158_add_4_1.INJECT1_0 = "NO";
    defparam sig_Vblank_158_add_4_1.INJECT1_1 = "NO";
    CCU2C sig_compt_front_Hsync_156_add_4_11 (.A0(sig_compt_front_Hsync[9]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(sig_compt_front_Hsync[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n1260), .COUT(n1261), 
          .S0(n76_adj_26), .S1(n75_adj_27));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156_add_4_11.INIT0 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_11.INIT1 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_11.INJECT1_0 = "NO";
    defparam sig_compt_front_Hsync_156_add_4_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut (.A(out_comp), .B(DE_c), .C(D_detect), .D(detect), 
         .Z(ODCK_c_enable_97)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B))) */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(173[9:35])
    defparam i1_4_lut_4_lut.init = 16'h4e44;
    LUT4 i1_2_lut_rep_7 (.A(Hsync_c), .B(DE_c), .Z(ODCK_c_enable_92)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_7.init = 16'heeee;
    LUT4 i11_4_lut (.A(sig_compt_front_Hsync[3]), .B(sig_compt_front_Hsync[11]), 
         .C(sig_compt_front_Hsync[13]), .D(sig_compt_front_Hsync[6]), .Z(n28_adj_65)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(sig_compt_front_Hsync[12]), .B(sig_compt_front_Hsync[8]), 
         .Z(n20)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i15_4_lut (.A(n17), .B(n30), .C(n26), .D(n18), .Z(out_comp_N_378)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i545_1_lut_rep_4_2_lut (.A(Hsync_c), .B(DE_c), .Z(ODCK_c_enable_17)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i545_1_lut_rep_4_2_lut.init = 16'h1111;
    LUT4 i1_2_lut (.A(sig_compt_front_Hsync[0]), .B(sig_compt_front_Hsync[10]), 
         .Z(n17)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(sig_compt_front_Hsync[14]), .B(sig_compt_front_Hsync[9]), 
         .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i12_4_lut (.A(sig_compt_front_Hsync[5]), .B(sig_compt_front_Hsync[7]), 
         .C(sig_compt_front_Hsync[2]), .D(sig_compt_front_Hsync[1]), .Z(n28)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut.init = 16'hfffe;
    CCU2C sig_Hdisp_cpt_147_add_4_17 (.A0(sig_Hdisp_cpt[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n1311), .S0(n70_adj_83));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147_add_4_17.INIT0 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_17.INIT1 = 16'h0000;
    defparam sig_Hdisp_cpt_147_add_4_17.INJECT1_0 = "NO";
    defparam sig_Hdisp_cpt_147_add_4_17.INJECT1_1 = "NO";
    CCU2C sig_Hdisp_cpt_147_add_4_15 (.A0(sig_Hdisp_cpt[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(sig_Hdisp_cpt[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n1310), .COUT(n1311), .S0(n72_adj_85), 
          .S1(n71_adj_84));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147_add_4_15.INIT0 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_15.INIT1 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_15.INJECT1_0 = "NO";
    defparam sig_Hdisp_cpt_147_add_4_15.INJECT1_1 = "NO";
    CCU2C sig_Hdisp_cpt_147_add_4_13 (.A0(sig_Hdisp_cpt[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(sig_Hdisp_cpt[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n1309), .COUT(n1310), .S0(n74_adj_87), 
          .S1(n73_adj_86));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147_add_4_13.INIT0 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_13.INIT1 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_13.INJECT1_0 = "NO";
    defparam sig_Hdisp_cpt_147_add_4_13.INJECT1_1 = "NO";
    CCU2C sig_Hdisp_cpt_147_add_4_11 (.A0(sig_Hdisp_cpt[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(sig_Hdisp_cpt[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n1308), .COUT(n1309), .S0(n76_adj_89), 
          .S1(n75_adj_88));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147_add_4_11.INIT0 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_11.INIT1 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_11.INJECT1_0 = "NO";
    defparam sig_Hdisp_cpt_147_add_4_11.INJECT1_1 = "NO";
    CCU2C sig_Hdisp_cpt_147_add_4_9 (.A0(sig_Hdisp_cpt[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(sig_Hdisp_cpt[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n1307), .COUT(n1308), .S0(n78_adj_91), 
          .S1(n77_adj_90));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147_add_4_9.INIT0 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_9.INIT1 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_9.INJECT1_0 = "NO";
    defparam sig_Hdisp_cpt_147_add_4_9.INJECT1_1 = "NO";
    CCU2C sig_Hsync_151_add_4_13 (.A0(Hsync_out_c_11), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hsync_out_c_12), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1293), .COUT(n1294), .S0(n74_adj_53), 
          .S1(n73_adj_52));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151_add_4_13.INIT0 = 16'haaa0;
    defparam sig_Hsync_151_add_4_13.INIT1 = 16'haaa0;
    defparam sig_Hsync_151_add_4_13.INJECT1_0 = "NO";
    defparam sig_Hsync_151_add_4_13.INJECT1_1 = "NO";
    CCU2C sig_Hsync_151_add_4_11 (.A0(Hsync_out_c_9), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hsync_out_c_10), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1292), .COUT(n1293), .S0(n76_adj_55), 
          .S1(n75_adj_54));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151_add_4_11.INIT0 = 16'haaa0;
    defparam sig_Hsync_151_add_4_11.INIT1 = 16'haaa0;
    defparam sig_Hsync_151_add_4_11.INJECT1_0 = "NO";
    defparam sig_Hsync_151_add_4_11.INJECT1_1 = "NO";
    CCU2C sig_Hblank_154_add_4_17 (.A0(Hblank_c_15), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n1279), .S0(n70_adj_16));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154_add_4_17.INIT0 = 16'haaa0;
    defparam sig_Hblank_154_add_4_17.INIT1 = 16'h0000;
    defparam sig_Hblank_154_add_4_17.INJECT1_0 = "NO";
    defparam sig_Hblank_154_add_4_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_2_lut_3_lut_1_lut (.A(DE_c), .Z(ODCK_c_enable_94)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_1_lut.init = 16'h5555;
    LUT4 Hsync_out_15__I_1_2_lut_rep_5 (.A(DE_c), .B(Hsync_c), .Z(n1380)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(107[7:31])
    defparam Hsync_out_15__I_1_2_lut_rep_5.init = 16'h4444;
    LUT4 i596_2_lut (.A(Vsync_c), .B(DE_c), .Z(ODCK_c_enable_95)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i596_2_lut.init = 16'h7777;
    LUT4 i497_1_lut (.A(Vsync_c), .Z(n1114)) /* synthesis lut_function=(!(A)) */ ;
    defparam i497_1_lut.init = 16'h5555;
    LUT4 i14_4_lut (.A(sig_compt_front_Hsync[10]), .B(n28_adj_65), .C(n20), 
         .D(sig_compt_front_Hsync[15]), .Z(n31)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i12_4_lut_adj_1 (.A(sig_compt_front_Hsync[4]), .B(sig_compt_front_Hsync[9]), 
         .C(sig_compt_front_Hsync[14]), .D(sig_compt_front_Hsync[5]), .Z(n29)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_1.init = 16'hfffe;
    LUT4 i2_2_lut (.A(sig_compt_front_Hsync[15]), .B(sig_compt_front_Hsync[12]), 
         .Z(n18)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1S3IX sig_Hblank_154__i16 (.D(n70_adj_16), .CK(ODCK_c), .CD(DE_c), 
            .Q(Hblank_c_15)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i16.GSR = "ENABLED";
    CCU2C sig_Hsync_151_add_4_9 (.A0(Hsync_out_c_7), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hsync_out_c_8), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1291), .COUT(n1292), .S0(n78_adj_57), 
          .S1(n77_adj_56));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151_add_4_9.INIT0 = 16'haaa0;
    defparam sig_Hsync_151_add_4_9.INIT1 = 16'haaa0;
    defparam sig_Hsync_151_add_4_9.INJECT1_0 = "NO";
    defparam sig_Hsync_151_add_4_9.INJECT1_1 = "NO";
    CCU2C sig_Hsync_151_add_4_7 (.A0(Hsync_out_c_5), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hsync_out_c_6), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1290), .COUT(n1291), .S0(n80_adj_59), 
          .S1(n79_adj_58));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151_add_4_7.INIT0 = 16'haaa0;
    defparam sig_Hsync_151_add_4_7.INIT1 = 16'haaa0;
    defparam sig_Hsync_151_add_4_7.INJECT1_0 = "NO";
    defparam sig_Hsync_151_add_4_7.INJECT1_1 = "NO";
    CCU2C sig_Hsync_151_add_4_5 (.A0(Hsync_out_c_3), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hsync_out_c_4), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1289), .COUT(n1290), .S0(n82_adj_61), 
          .S1(n81_adj_60));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151_add_4_5.INIT0 = 16'haaa0;
    defparam sig_Hsync_151_add_4_5.INIT1 = 16'haaa0;
    defparam sig_Hsync_151_add_4_5.INJECT1_0 = "NO";
    defparam sig_Hsync_151_add_4_5.INJECT1_1 = "NO";
    CCU2C sig_Hsync_151_add_4_3 (.A0(Hsync_out_c_1), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Hsync_out_c_2), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1288), .COUT(n1289), .S0(n84_adj_63), 
          .S1(n83_adj_62));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151_add_4_3.INIT0 = 16'haaa0;
    defparam sig_Hsync_151_add_4_3.INIT1 = 16'haaa0;
    defparam sig_Hsync_151_add_4_3.INJECT1_0 = "NO";
    defparam sig_Hsync_151_add_4_3.INJECT1_1 = "NO";
    CCU2C sig_Hsync_151_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Hsync_out_c_0), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n1288), .S1(n85_adj_64));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151_add_4_1.INIT0 = 16'h0000;
    defparam sig_Hsync_151_add_4_1.INIT1 = 16'h555f;
    defparam sig_Hsync_151_add_4_1.INJECT1_0 = "NO";
    defparam sig_Hsync_151_add_4_1.INJECT1_1 = "NO";
    CCU2C sig_Vsync_153_add_4_17 (.A0(Vsync_out_c_15), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n1287), .S0(n70_adj_33));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153_add_4_17.INIT0 = 16'haaa0;
    defparam sig_Vsync_153_add_4_17.INIT1 = 16'h0000;
    defparam sig_Vsync_153_add_4_17.INJECT1_0 = "NO";
    defparam sig_Vsync_153_add_4_17.INJECT1_1 = "NO";
    CCU2C sig_Vsync_153_add_4_15 (.A0(Vsync_out_c_13), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vsync_out_c_14), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1286), .COUT(n1287), .S0(n72_adj_35), 
          .S1(n71_adj_34));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153_add_4_15.INIT0 = 16'haaa0;
    defparam sig_Vsync_153_add_4_15.INIT1 = 16'haaa0;
    defparam sig_Vsync_153_add_4_15.INJECT1_0 = "NO";
    defparam sig_Vsync_153_add_4_15.INJECT1_1 = "NO";
    CCU2C sig_Vsync_153_add_4_13 (.A0(Vsync_out_c_11), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vsync_out_c_12), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1285), .COUT(n1286), .S0(n74_adj_37), 
          .S1(n73_adj_36));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153_add_4_13.INIT0 = 16'haaa0;
    defparam sig_Vsync_153_add_4_13.INIT1 = 16'haaa0;
    defparam sig_Vsync_153_add_4_13.INJECT1_0 = "NO";
    defparam sig_Vsync_153_add_4_13.INJECT1_1 = "NO";
    CCU2C sig_Vsync_153_add_4_11 (.A0(Vsync_out_c_9), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vsync_out_c_10), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1284), .COUT(n1285), .S0(n76_adj_39), 
          .S1(n75_adj_38));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153_add_4_11.INIT0 = 16'haaa0;
    defparam sig_Vsync_153_add_4_11.INIT1 = 16'haaa0;
    defparam sig_Vsync_153_add_4_11.INJECT1_0 = "NO";
    defparam sig_Vsync_153_add_4_11.INJECT1_1 = "NO";
    CCU2C sig_Vsync_153_add_4_9 (.A0(Vsync_out_c_7), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vsync_out_c_8), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1283), .COUT(n1284), .S0(n78_adj_41), 
          .S1(n77_adj_40));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153_add_4_9.INIT0 = 16'haaa0;
    defparam sig_Vsync_153_add_4_9.INIT1 = 16'haaa0;
    defparam sig_Vsync_153_add_4_9.INJECT1_0 = "NO";
    defparam sig_Vsync_153_add_4_9.INJECT1_1 = "NO";
    CCU2C sig_Vsync_153_add_4_7 (.A0(Vsync_out_c_5), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vsync_out_c_6), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1282), .COUT(n1283), .S0(n80_adj_43), 
          .S1(n79_adj_42));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153_add_4_7.INIT0 = 16'haaa0;
    defparam sig_Vsync_153_add_4_7.INIT1 = 16'haaa0;
    defparam sig_Vsync_153_add_4_7.INJECT1_0 = "NO";
    defparam sig_Vsync_153_add_4_7.INJECT1_1 = "NO";
    CCU2C sig_Vsync_153_add_4_5 (.A0(Vsync_out_c_3), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vsync_out_c_4), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1281), .COUT(n1282), .S0(n82_adj_45), 
          .S1(n81_adj_44));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153_add_4_5.INIT0 = 16'haaa0;
    defparam sig_Vsync_153_add_4_5.INIT1 = 16'haaa0;
    defparam sig_Vsync_153_add_4_5.INJECT1_0 = "NO";
    defparam sig_Vsync_153_add_4_5.INJECT1_1 = "NO";
    CCU2C sig_Vsync_153_add_4_3 (.A0(Vsync_out_c_1), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vsync_out_c_2), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1280), .COUT(n1281), .S0(n84_adj_47), 
          .S1(n83_adj_46));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153_add_4_3.INIT0 = 16'haaa0;
    defparam sig_Vsync_153_add_4_3.INIT1 = 16'haaa0;
    defparam sig_Vsync_153_add_4_3.INJECT1_0 = "NO";
    defparam sig_Vsync_153_add_4_3.INJECT1_1 = "NO";
    CCU2C sig_Vsync_153_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Vsync_out_c_0), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n1280), .S1(n85_adj_48));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153_add_4_1.INIT0 = 16'h0000;
    defparam sig_Vsync_153_add_4_1.INIT1 = 16'h555f;
    defparam sig_Vsync_153_add_4_1.INJECT1_0 = "NO";
    defparam sig_Vsync_153_add_4_1.INJECT1_1 = "NO";
    CCU2C sig_Hdisp_cpt_147_add_4_5 (.A0(sig_Hdisp_cpt[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(sig_Hdisp_cpt[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n1305), .COUT(n1306), .S0(n82_adj_95), 
          .S1(n81_adj_94));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147_add_4_5.INIT0 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_5.INIT1 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_5.INJECT1_0 = "NO";
    defparam sig_Hdisp_cpt_147_add_4_5.INJECT1_1 = "NO";
    FD1S3IX sig_Hblank_154__i15 (.D(n71_adj_15), .CK(ODCK_c), .CD(DE_c), 
            .Q(Hblank_c_14)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i15.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i14 (.D(n72_adj_14), .CK(ODCK_c), .CD(DE_c), 
            .Q(Hblank_c_13)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i14.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i13 (.D(n73), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_12)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i13.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i12 (.D(n74), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_11)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i12.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i11 (.D(n75), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_10)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i11.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i10 (.D(n76), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_9)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i10.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i9 (.D(n77), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_8)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i9.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i8 (.D(n78), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_7)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i8.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i7 (.D(n79), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_6)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i7.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i6 (.D(n80), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_5)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i6.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i5 (.D(n81), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_4)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i5.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i4 (.D(n82), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_3)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i4.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i3 (.D(n83), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_2)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i3.GSR = "ENABLED";
    FD1S3IX sig_Hblank_154__i2 (.D(n84), .CK(ODCK_c), .CD(DE_c), .Q(Hblank_c_1)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hblank_154__i2.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i16 (.D(sig_Hdisp_cpt[15]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_15)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i16.GSR = "ENABLED";
    CCU2C sig_Hdisp_cpt_147_add_4_3 (.A0(sig_Hdisp_cpt[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(sig_Hdisp_cpt[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n1304), .COUT(n1305), .S0(n84_adj_97), 
          .S1(n83_adj_96));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147_add_4_3.INIT0 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_3.INIT1 = 16'haaa0;
    defparam sig_Hdisp_cpt_147_add_4_3.INJECT1_0 = "NO";
    defparam sig_Hdisp_cpt_147_add_4_3.INJECT1_1 = "NO";
    CCU2C sig_Hdisp_cpt_147_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(sig_Hdisp_cpt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n1304), .S1(n85_adj_98));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147_add_4_1.INIT0 = 16'h0000;
    defparam sig_Hdisp_cpt_147_add_4_1.INIT1 = 16'h555f;
    defparam sig_Hdisp_cpt_147_add_4_1.INJECT1_0 = "NO";
    defparam sig_Hdisp_cpt_147_add_4_1.INJECT1_1 = "NO";
    CCU2C sig_Vdisp_149_add_4_17 (.A0(Vdisp_c_15), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n1303), .S0(n70_adj_67));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149_add_4_17.INIT0 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_17.INIT1 = 16'h0000;
    defparam sig_Vdisp_149_add_4_17.INJECT1_0 = "NO";
    defparam sig_Vdisp_149_add_4_17.INJECT1_1 = "NO";
    CCU2C sig_Vdisp_149_add_4_15 (.A0(Vdisp_c_13), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vdisp_c_14), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1302), .COUT(n1303), .S0(n72_adj_69), 
          .S1(n71_adj_68));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149_add_4_15.INIT0 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_15.INIT1 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_15.INJECT1_0 = "NO";
    defparam sig_Vdisp_149_add_4_15.INJECT1_1 = "NO";
    CCU2C sig_Vdisp_149_add_4_13 (.A0(Vdisp_c_11), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vdisp_c_12), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1301), .COUT(n1302), .S0(n74_adj_71), 
          .S1(n73_adj_70));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149_add_4_13.INIT0 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_13.INIT1 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_13.INJECT1_0 = "NO";
    defparam sig_Vdisp_149_add_4_13.INJECT1_1 = "NO";
    CCU2C sig_Vdisp_149_add_4_11 (.A0(Vdisp_c_9), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vdisp_c_10), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1300), .COUT(n1301), .S0(n76_adj_73), 
          .S1(n75_adj_72));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149_add_4_11.INIT0 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_11.INIT1 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_11.INJECT1_0 = "NO";
    defparam sig_Vdisp_149_add_4_11.INJECT1_1 = "NO";
    CCU2C sig_Vdisp_149_add_4_9 (.A0(Vdisp_c_7), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vdisp_c_8), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1299), .COUT(n1300), .S0(n78_adj_75), 
          .S1(n77_adj_74));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149_add_4_9.INIT0 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_9.INIT1 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_9.INJECT1_0 = "NO";
    defparam sig_Vdisp_149_add_4_9.INJECT1_1 = "NO";
    CCU2C sig_Vdisp_149_add_4_7 (.A0(Vdisp_c_5), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vdisp_c_6), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1298), .COUT(n1299), .S0(n80_adj_77), 
          .S1(n79_adj_76));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149_add_4_7.INIT0 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_7.INIT1 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_7.INJECT1_0 = "NO";
    defparam sig_Vdisp_149_add_4_7.INJECT1_1 = "NO";
    CCU2C sig_Vdisp_149_add_4_5 (.A0(Vdisp_c_3), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vdisp_c_4), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1297), .COUT(n1298), .S0(n82_adj_79), 
          .S1(n81_adj_78));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149_add_4_5.INIT0 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_5.INIT1 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_5.INJECT1_0 = "NO";
    defparam sig_Vdisp_149_add_4_5.INJECT1_1 = "NO";
    CCU2C sig_Vdisp_149_add_4_3 (.A0(Vdisp_c_1), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(Vdisp_c_2), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n1296), .COUT(n1297), .S0(n84_adj_81), 
          .S1(n83_adj_80));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149_add_4_3.INIT0 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_3.INIT1 = 16'haaa0;
    defparam sig_Vdisp_149_add_4_3.INJECT1_0 = "NO";
    defparam sig_Vdisp_149_add_4_3.INJECT1_1 = "NO";
    CCU2C sig_Vdisp_149_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Vdisp_c_0), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n1296), .S1(n85_adj_82));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149_add_4_1.INIT0 = 16'h0000;
    defparam sig_Vdisp_149_add_4_1.INIT1 = 16'h555f;
    defparam sig_Vdisp_149_add_4_1.INJECT1_0 = "NO";
    defparam sig_Vdisp_149_add_4_1.INJECT1_1 = "NO";
    CCU2C sig_compt_front_Hsync_156_add_4_9 (.A0(sig_compt_front_Hsync[7]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(sig_compt_front_Hsync[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n1259), .COUT(n1260), 
          .S0(n78_adj_24), .S1(n77_adj_25));   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156_add_4_9.INIT0 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_9.INIT1 = 16'haaa0;
    defparam sig_compt_front_Hsync_156_add_4_9.INJECT1_0 = "NO";
    defparam sig_compt_front_Hsync_156_add_4_9.INJECT1_1 = "NO";
    FD1P3IX sig_Vblank_158__i2 (.D(n84_adj_2), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_1)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i2.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i15 (.D(sig_Hdisp_cpt[14]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_14)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i15.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i14 (.D(sig_Hdisp_cpt[13]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_13)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i14.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i13 (.D(sig_Hdisp_cpt[12]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_12)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i13.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i12 (.D(sig_Hdisp_cpt[11]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_11)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i12.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i11 (.D(sig_Hdisp_cpt[10]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_10)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i11.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i10 (.D(sig_Hdisp_cpt[9]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_9)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i10.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i9 (.D(sig_Hdisp_cpt[8]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_8)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i9.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i8 (.D(sig_Hdisp_cpt[7]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_7)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i8.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i7 (.D(sig_Hdisp_cpt[6]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_6)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i7.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i6 (.D(sig_Hdisp_cpt[5]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_5)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i6.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i5 (.D(sig_Hdisp_cpt[4]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_4)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i5.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i4 (.D(sig_Hdisp_cpt[3]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_3)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i4.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i3 (.D(sig_Hdisp_cpt[2]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_2)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i3.GSR = "ENABLED";
    FD1P3AX sig_Hdisp_i0_i2 (.D(sig_Hdisp_cpt[1]), .SP(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hdisp_c_1)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(77[1] 86[9])
    defparam sig_Hdisp_i0_i2.GSR = "ENABLED";
    LUT4 i10_4_lut (.A(sig_compt_front_Hsync[8]), .B(sig_compt_front_Hsync[13]), 
         .C(sig_compt_front_Hsync[3]), .D(sig_compt_front_Hsync[11]), .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut.init = 16'hfffe;
    FD1P3IX sig_Vblank_158__i3 (.D(n83_adj_3), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_2)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i3.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i4 (.D(n82_adj_4), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_3)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i4.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i5 (.D(n81_adj_5), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_4)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i5.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i6 (.D(n80_adj_6), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_5)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i6.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i7 (.D(n79_adj_7), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_6)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i7.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i8 (.D(n78_adj_8), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_7)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i8.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i9 (.D(n77_adj_9), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_8)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i9.GSR = "ENABLED";
    LUT4 i412_2_lut_3_lut_4_lut (.A(DE_c), .B(Vsync_c), .C(detect_DE), 
         .D(D_detect_DE), .Z(n1084)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(39[1:3])
    defparam i412_2_lut_3_lut_4_lut.init = 16'h4044;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VLO i1 (.Z(GND_net));
    LUT4 i16_4_lut (.A(n31), .B(n29), .C(n25), .D(n26_adj_66), .Z(ODCK_c_enable_96)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16_4_lut.init = 16'hfffe;
    FD1P3IX sig_compt_front_Hsync_156__i15 (.D(n70_adj_32), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[15])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i15.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i10 (.D(n76_adj_10), .SP(ODCK_c_enable_97), 
            .CD(n1381), .CK(ODCK_c), .Q(Vblank_c_9)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i10.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i11 (.D(n75_adj_11), .SP(ODCK_c_enable_97), 
            .CD(n1381), .CK(ODCK_c), .Q(Vblank_c_10)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i11.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i12 (.D(n74_adj_12), .SP(ODCK_c_enable_97), 
            .CD(n1381), .CK(ODCK_c), .Q(Vblank_c_11)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i12.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i13 (.D(n73_adj_13), .SP(ODCK_c_enable_97), 
            .CD(n1381), .CK(ODCK_c), .Q(Vblank_c_12)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i13.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i14 (.D(n72), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_13)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i14.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i15 (.D(n71), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_14)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i15.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i16 (.D(n70), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_15)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i16.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i2 (.D(n84_adj_47), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_1)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i2.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i3 (.D(n83_adj_46), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_2)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i3.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i4 (.D(n82_adj_45), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_3)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i4.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i5 (.D(n81_adj_44), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_4)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i5.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i6 (.D(n80_adj_43), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_5)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i6.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i7 (.D(n79_adj_42), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_6)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i7.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i8 (.D(n78_adj_41), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_7)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i8.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i9 (.D(n77_adj_40), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_8)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i9.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i10 (.D(n76_adj_39), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_9)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i10.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i11 (.D(n75_adj_38), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_10)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i11.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i12 (.D(n74_adj_37), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_11)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i12.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i13 (.D(n73_adj_36), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_12)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i13.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i14 (.D(n72_adj_35), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_13)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i14.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i15 (.D(n71_adj_34), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_14)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i15.GSR = "ENABLED";
    FD1P3IX sig_Vsync_153__i16 (.D(n70_adj_33), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_15)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i16.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i2 (.D(n84_adj_63), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_1)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i2.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i3 (.D(n83_adj_62), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_2)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i3.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i4 (.D(n82_adj_61), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_3)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i4.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i5 (.D(n81_adj_60), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_4)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i5.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i6 (.D(n80_adj_59), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_5)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i6.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i7 (.D(n79_adj_58), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_6)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i7.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i8 (.D(n78_adj_57), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_7)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i8.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i9 (.D(n77_adj_56), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_8)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i9.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i10 (.D(n76_adj_55), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_9)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i10.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i11 (.D(n75_adj_54), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_10)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i11.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i12 (.D(n74_adj_53), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_11)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i12.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i13 (.D(n73_adj_52), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_12)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i13.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i14 (.D(n72_adj_51), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_13)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i14.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i15 (.D(n71_adj_50), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_14)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i15.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i16 (.D(n70_adj_49), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_15)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i16.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i2 (.D(n84_adj_81), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_1)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i2.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i3 (.D(n83_adj_80), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_2)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i3.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i4 (.D(n82_adj_79), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_3)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i4.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i5 (.D(n81_adj_78), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_4)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i5.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i6 (.D(n80_adj_77), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_5)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i6.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i7 (.D(n79_adj_76), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_6)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i7.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i8 (.D(n78_adj_75), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_7)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i8.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i9 (.D(n77_adj_74), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_8)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i9.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i10 (.D(n76_adj_73), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_9)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i10.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i11 (.D(n75_adj_72), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_10)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i11.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i12 (.D(n74_adj_71), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_11)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i12.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i13 (.D(n73_adj_70), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_12)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i13.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i14 (.D(n72_adj_69), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_13)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i14.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i15 (.D(n71_adj_68), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_14)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i15.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i16 (.D(n70_adj_67), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_15)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i16.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i14 (.D(n71_adj_31), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[14])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i14.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i13 (.D(n72_adj_30), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[13])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i13.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i12 (.D(n73_adj_29), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[12])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i12.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i11 (.D(n74_adj_28), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[11])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i11.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i10 (.D(n75_adj_27), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[10])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i10.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i9 (.D(n76_adj_26), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i9.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i8 (.D(n77_adj_25), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i8.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i7 (.D(n78_adj_24), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i7.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i6 (.D(n79_adj_23), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i6.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i5 (.D(n80_adj_22), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i5.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i4 (.D(n81_adj_21), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i4.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i3 (.D(n82_adj_20), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i3.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i2 (.D(n83_adj_19), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i2.GSR = "ENABLED";
    FD1P3IX sig_compt_front_Hsync_156__i1 (.D(n84_adj_18), .SP(rising_Hsync), 
            .CD(DE_c), .CK(ODCK_c), .Q(sig_compt_front_Hsync[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_compt_front_Hsync_156__i1.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i1 (.D(n84_adj_97), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i1.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i2 (.D(n83_adj_96), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i2.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i3 (.D(n82_adj_95), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i3.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i4 (.D(n81_adj_94), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i4.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i5 (.D(n80_adj_93), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i5.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i6 (.D(n79_adj_92), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i6.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i7 (.D(n78_adj_91), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i7.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i8 (.D(n77_adj_90), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i8.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i9 (.D(n76_adj_89), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i9.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i10 (.D(n75_adj_88), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i10.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i11 (.D(n74_adj_87), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i11.GSR = "ENABLED";
    OB Hdisp_pad_7 (.I(Hdisp_c_7), .O(Hdisp[7]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    OB Hdisp_pad_6 (.I(Hdisp_c_6), .O(Hdisp[6]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    OB Hdisp_pad_5 (.I(Hdisp_c_5), .O(Hdisp[5]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    OB Hdisp_pad_4 (.I(Hdisp_c_4), .O(Hdisp[4]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    OB Hdisp_pad_3 (.I(Hdisp_c_3), .O(Hdisp[3]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    OB Hdisp_pad_2 (.I(Hdisp_c_2), .O(Hdisp[2]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    OB Hdisp_pad_1 (.I(Hdisp_c_1), .O(Hdisp[1]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    OB Hdisp_pad_0 (.I(Hdisp_c_0), .O(Hdisp[0]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(44[1:6])
    OB Vdisp_pad_15 (.I(Vdisp_c_15), .O(Vdisp[15]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_14 (.I(Vdisp_c_14), .O(Vdisp[14]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_13 (.I(Vdisp_c_13), .O(Vdisp[13]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_12 (.I(Vdisp_c_12), .O(Vdisp[12]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_11 (.I(Vdisp_c_11), .O(Vdisp[11]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_10 (.I(Vdisp_c_10), .O(Vdisp[10]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_9 (.I(Vdisp_c_9), .O(Vdisp[9]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_8 (.I(Vdisp_c_8), .O(Vdisp[8]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_7 (.I(Vdisp_c_7), .O(Vdisp[7]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_6 (.I(Vdisp_c_6), .O(Vdisp[6]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_5 (.I(Vdisp_c_5), .O(Vdisp[5]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_4 (.I(Vdisp_c_4), .O(Vdisp[4]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_3 (.I(Vdisp_c_3), .O(Vdisp[3]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_2 (.I(Vdisp_c_2), .O(Vdisp[2]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_1 (.I(Vdisp_c_1), .O(Vdisp[1]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Vdisp_pad_0 (.I(Vdisp_c_0), .O(Vdisp[0]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(45[1:6])
    OB Hblank_pad_15 (.I(Hblank_c_15), .O(Hblank[15]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_14 (.I(Hblank_c_14), .O(Hblank[14]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_13 (.I(Hblank_c_13), .O(Hblank[13]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_12 (.I(Hblank_c_12), .O(Hblank[12]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_11 (.I(Hblank_c_11), .O(Hblank[11]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_10 (.I(Hblank_c_10), .O(Hblank[10]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_9 (.I(Hblank_c_9), .O(Hblank[9]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_8 (.I(Hblank_c_8), .O(Hblank[8]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_7 (.I(Hblank_c_7), .O(Hblank[7]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_6 (.I(Hblank_c_6), .O(Hblank[6]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_5 (.I(Hblank_c_5), .O(Hblank[5]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_4 (.I(Hblank_c_4), .O(Hblank[4]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_3 (.I(Hblank_c_3), .O(Hblank[3]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_2 (.I(Hblank_c_2), .O(Hblank[2]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_1 (.I(Hblank_c_1), .O(Hblank[1]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Hblank_pad_0 (.I(Hblank_c_0), .O(Hblank[0]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(46[1:7])
    OB Vblank_pad_15 (.I(Vblank_c_15), .O(Vblank[15]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_14 (.I(Vblank_c_14), .O(Vblank[14]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_13 (.I(Vblank_c_13), .O(Vblank[13]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_12 (.I(Vblank_c_12), .O(Vblank[12]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_11 (.I(Vblank_c_11), .O(Vblank[11]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_10 (.I(Vblank_c_10), .O(Vblank[10]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_9 (.I(Vblank_c_9), .O(Vblank[9]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_8 (.I(Vblank_c_8), .O(Vblank[8]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_7 (.I(Vblank_c_7), .O(Vblank[7]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_6 (.I(Vblank_c_6), .O(Vblank[6]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_5 (.I(Vblank_c_5), .O(Vblank[5]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_4 (.I(Vblank_c_4), .O(Vblank[4]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_3 (.I(Vblank_c_3), .O(Vblank[3]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_2 (.I(Vblank_c_2), .O(Vblank[2]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_1 (.I(Vblank_c_1), .O(Vblank[1]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Vblank_pad_0 (.I(Vblank_c_0), .O(Vblank[0]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(47[1:7])
    OB Hsync_out_pad_15 (.I(Hsync_out_c_15), .O(Hsync_out[15]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_14 (.I(Hsync_out_c_14), .O(Hsync_out[14]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_13 (.I(Hsync_out_c_13), .O(Hsync_out[13]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_12 (.I(Hsync_out_c_12), .O(Hsync_out[12]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_11 (.I(Hsync_out_c_11), .O(Hsync_out[11]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_10 (.I(Hsync_out_c_10), .O(Hsync_out[10]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_9 (.I(Hsync_out_c_9), .O(Hsync_out[9]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_8 (.I(Hsync_out_c_8), .O(Hsync_out[8]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_7 (.I(Hsync_out_c_7), .O(Hsync_out[7]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_6 (.I(Hsync_out_c_6), .O(Hsync_out[6]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_5 (.I(Hsync_out_c_5), .O(Hsync_out[5]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_4 (.I(Hsync_out_c_4), .O(Hsync_out[4]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_3 (.I(Hsync_out_c_3), .O(Hsync_out[3]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_2 (.I(Hsync_out_c_2), .O(Hsync_out[2]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_1 (.I(Hsync_out_c_1), .O(Hsync_out[1]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Hsync_out_pad_0 (.I(Hsync_out_c_0), .O(Hsync_out[0]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(48[1:10])
    OB Vsync_out_pad_15 (.I(Vsync_out_c_15), .O(Vsync_out[15]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_14 (.I(Vsync_out_c_14), .O(Vsync_out[14]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_13 (.I(Vsync_out_c_13), .O(Vsync_out[13]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_12 (.I(Vsync_out_c_12), .O(Vsync_out[12]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_11 (.I(Vsync_out_c_11), .O(Vsync_out[11]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_10 (.I(Vsync_out_c_10), .O(Vsync_out[10]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_9 (.I(Vsync_out_c_9), .O(Vsync_out[9]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_8 (.I(Vsync_out_c_8), .O(Vsync_out[8]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_7 (.I(Vsync_out_c_7), .O(Vsync_out[7]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_6 (.I(Vsync_out_c_6), .O(Vsync_out[6]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_5 (.I(Vsync_out_c_5), .O(Vsync_out[5]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_4 (.I(Vsync_out_c_4), .O(Vsync_out[4]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_3 (.I(Vsync_out_c_3), .O(Vsync_out[3]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_2 (.I(Vsync_out_c_2), .O(Vsync_out[2]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_1 (.I(Vsync_out_c_1), .O(Vsync_out[1]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    OB Vsync_out_pad_0 (.I(Vsync_out_c_0), .O(Vsync_out[0]));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(49[1:10])
    IB DE_pad (.I(DE), .O(DE_c));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(39[1:3])
    IB Vsync_pad (.I(Vsync), .O(Vsync_c));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(40[1:6])
    IB Hsync_pad (.I(Hsync), .O(Hsync_c));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(41[1:6])
    IB ODCK_pad (.I(ODCK), .O(ODCK_c));   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(42[1:5])
    FD1P3IX sig_Hdisp_cpt_147__i12 (.D(n73_adj_86), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i12.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i13 (.D(n72_adj_85), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i13.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i14 (.D(n71_adj_84), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[14])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i14.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i15 (.D(n70_adj_83), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[15])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i15.GSR = "ENABLED";
    FD1P3IX sig_Hdisp_cpt_147__i0 (.D(n85_adj_98), .SP(ODCK_c_enable_92), 
            .CD(n1380), .CK(ODCK_c), .Q(sig_Hdisp_cpt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hdisp_cpt_147__i0.GSR = "ENABLED";
    FD1P3IX sig_Vdisp_149__i1 (.D(n85_adj_82), .SP(ODCK_c_enable_93), .CD(n1084), 
            .CK(ODCK_c), .Q(Vdisp_c_0)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vdisp_149__i1.GSR = "ENABLED";
    FD1P3IX sig_Hsync_151__i1 (.D(n85_adj_64), .SP(ODCK_c_enable_94), .CD(ODCK_c_enable_17), 
            .CK(ODCK_c), .Q(Hsync_out_c_0)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Hsync_151__i1.GSR = "ENABLED";
    LUT4 rising_Hsync_I_0_2_lut (.A(D_detect), .B(detect), .Z(rising_Hsync)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(187[5:36])
    defparam rising_Hsync_I_0_2_lut.init = 16'h4444;
    FD1P3IX sig_Vsync_153__i1 (.D(n85_adj_48), .SP(ODCK_c_enable_95), .CD(n1114), 
            .CK(ODCK_c), .Q(Vsync_out_c_0)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vsync_153__i1.GSR = "ENABLED";
    LUT4 i14_4_lut_adj_2 (.A(sig_compt_front_Hsync[6]), .B(n28), .C(n22), 
         .D(sig_compt_front_Hsync[4]), .Z(n30)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut_adj_2.init = 16'hfffe;
    FD1P3IX out_comp_89 (.D(out_comp_N_378), .SP(ODCK_c_enable_96), .CD(DE_c), 
            .CK(ODCK_c), .Q(out_comp)) /* synthesis lse_init_val=0 */ ;   // /home/diamond/SharedFolder/DiamondProjFolder/test_DVI.vhd(158[1] 164[9])
    defparam out_comp_89.GSR = "ENABLED";
    FD1P3IX sig_Vblank_158__i1 (.D(n85_adj_1), .SP(ODCK_c_enable_97), .CD(n1381), 
            .CK(ODCK_c), .Q(Vblank_c_0)) /* synthesis syn_use_carry_chain=1 */ ;   // /usr/local/diamond/3.11_x64/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam sig_Vblank_158__i1.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.3.469 */
/* Module Version: 6.5 */
/* /usr/local/diamond/3.11_x64/ispfpga/bin/lin64/scuba -w -bus_exp 7 -bb -arch ep5c00 -type bram -wp 10 -rp 0011 -data_width 1 -num_rows 2 -rdata_width 1 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpEbnonesadr112112115216de -pmi -lang verilog  */
/* Mon Mar 29 18:50:34 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpEbnonesadr112112115216de (WrAddress, RdAddress, Data, 
    WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [0:0] WrAddress;
    input wire [0:0] RdAddress;
    input wire [0:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [0:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpEbnonesadr112112115216de_0_0_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr112112115216de_0_0_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr112112115216de_0_0_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr112112115216de_0_0_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr112112115216de_0_0_0.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr112112115216de_0_0_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr112112115216de_0_0_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr112112115216de_0_0_0.DATA_WIDTH_B = 1 ;
    defparam pmi_ram_dpEbnonesadr112112115216de_0_0_0.DATA_WIDTH_A = 1 ;
    DP16KC pmi_ram_dpEbnonesadr112112115216de_0_0_0 (.DIA0(scuba_vlo), .DIA1(scuba_vlo), 
        .DIA2(scuba_vlo), .DIA3(scuba_vlo), .DIA4(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA6(scuba_vlo), .DIA7(scuba_vlo), .DIA8(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA10(scuba_vlo), .DIA11(Data[0]), .DIA12(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), .DIA17(scuba_vlo), 
        .ADA0(WrAddress[0]), .ADA1(scuba_vlo), .ADA2(scuba_vlo), .ADA3(scuba_vlo), 
        .ADA4(scuba_vlo), .ADA5(scuba_vlo), .ADA6(scuba_vlo), .ADA7(scuba_vlo), 
        .ADA8(scuba_vlo), .ADA9(scuba_vlo), .ADA10(scuba_vlo), .ADA11(scuba_vlo), 
        .ADA12(scuba_vlo), .ADA13(scuba_vlo), .CEA(WrClockEn), .CLKA(WrClock), 
        .OCEA(WrClockEn), .WEA(WE), .CSA0(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA2(scuba_vlo), .RSTA(Reset), .DIB0(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), .DIB17(scuba_vlo), 
        .ADB0(RdAddress[0]), .ADB1(scuba_vlo), .ADB2(scuba_vlo), .ADB3(scuba_vlo), 
        .ADB4(scuba_vlo), .ADB5(scuba_vlo), .ADB6(scuba_vlo), .ADB7(scuba_vlo), 
        .ADB8(scuba_vlo), .ADB9(scuba_vlo), .ADB10(scuba_vlo), .ADB11(scuba_vlo), 
        .ADB12(scuba_vlo), .ADB13(scuba_vlo), .CEB(RdClockEn), .CLKB(RdClock), 
        .OCEB(RdClockEn), .WEB(scuba_vlo), .CSB0(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB2(scuba_vlo), .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), 
        .DOA4(), .DOA5(), .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), 
        .DOA11(), .DOA12(), .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), 
        .DOB0(Q[0]), .DOB1(), .DOB2(), .DOB3(), .DOB4(), .DOB5(), .DOB6(), 
        .DOB7(), .DOB8(), .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), 
        .DOB14(), .DOB15(), .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr112112115216de__PMIP__2__1__1B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpEbnonesadr112112115216de_0_0_0 MEM_LPC_FILE pmi_ram_dpEbnonesadr112112115216de__PMIP__2__1__1B
    // exemplar attribute pmi_ram_dpEbnonesadr112112115216de_0_0_0 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr112112115216de_0_0_0 RESETMODE SYNC
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.3.469 */
/* Module Version: 6.5 */
/* /usr/local/diamond/3.11_x64/ispfpga/bin/lin64/scuba -w -bus_exp 7 -bb -arch ep5c00 -type bram -wp 10 -rp 0011 -data_width 99 -num_rows 16384 -rdata_width 99 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpEbnonesadr991416384991416384122adcc5 -pmi -lang verilog  */
/* Mon Mar 29 18:50:33 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpEbnonesadr991416384991416384122adcc5 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [13:0] WrAddress;
    input wire [13:0] RdAddress;
    input wire [98:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [98:0] Q;

    wire scuba_vhi;
    wire raddr11_ff;
    wire raddr12_ff;
    wire scuba_vlo;
    wire raddr13_ff;
    wire mdout1_7_0;
    wire mdout1_6_0;
    wire mdout1_5_0;
    wire mdout1_4_0;
    wire mdout1_3_0;
    wire mdout1_2_0;
    wire mdout1_1_0;
    wire mdout1_0_0;
    wire mdout1_7_1;
    wire mdout1_6_1;
    wire mdout1_5_1;
    wire mdout1_4_1;
    wire mdout1_3_1;
    wire mdout1_2_1;
    wire mdout1_1_1;
    wire mdout1_0_1;
    wire mdout1_7_2;
    wire mdout1_6_2;
    wire mdout1_5_2;
    wire mdout1_4_2;
    wire mdout1_3_2;
    wire mdout1_2_2;
    wire mdout1_1_2;
    wire mdout1_0_2;
    wire mdout1_7_3;
    wire mdout1_6_3;
    wire mdout1_5_3;
    wire mdout1_4_3;
    wire mdout1_3_3;
    wire mdout1_2_3;
    wire mdout1_1_3;
    wire mdout1_0_3;
    wire mdout1_7_4;
    wire mdout1_6_4;
    wire mdout1_5_4;
    wire mdout1_4_4;
    wire mdout1_3_4;
    wire mdout1_2_4;
    wire mdout1_1_4;
    wire mdout1_0_4;
    wire mdout1_7_5;
    wire mdout1_6_5;
    wire mdout1_5_5;
    wire mdout1_4_5;
    wire mdout1_3_5;
    wire mdout1_2_5;
    wire mdout1_1_5;
    wire mdout1_0_5;
    wire mdout1_7_6;
    wire mdout1_6_6;
    wire mdout1_5_6;
    wire mdout1_4_6;
    wire mdout1_3_6;
    wire mdout1_2_6;
    wire mdout1_1_6;
    wire mdout1_0_6;
    wire mdout1_7_7;
    wire mdout1_6_7;
    wire mdout1_5_7;
    wire mdout1_4_7;
    wire mdout1_3_7;
    wire mdout1_2_7;
    wire mdout1_1_7;
    wire mdout1_0_7;
    wire mdout1_7_8;
    wire mdout1_6_8;
    wire mdout1_5_8;
    wire mdout1_4_8;
    wire mdout1_3_8;
    wire mdout1_2_8;
    wire mdout1_1_8;
    wire mdout1_0_8;
    wire mdout1_7_9;
    wire mdout1_6_9;
    wire mdout1_5_9;
    wire mdout1_4_9;
    wire mdout1_3_9;
    wire mdout1_2_9;
    wire mdout1_1_9;
    wire mdout1_0_9;
    wire mdout1_7_10;
    wire mdout1_6_10;
    wire mdout1_5_10;
    wire mdout1_4_10;
    wire mdout1_3_10;
    wire mdout1_2_10;
    wire mdout1_1_10;
    wire mdout1_0_10;
    wire mdout1_7_11;
    wire mdout1_6_11;
    wire mdout1_5_11;
    wire mdout1_4_11;
    wire mdout1_3_11;
    wire mdout1_2_11;
    wire mdout1_1_11;
    wire mdout1_0_11;
    wire mdout1_7_12;
    wire mdout1_6_12;
    wire mdout1_5_12;
    wire mdout1_4_12;
    wire mdout1_3_12;
    wire mdout1_2_12;
    wire mdout1_1_12;
    wire mdout1_0_12;
    wire mdout1_7_13;
    wire mdout1_6_13;
    wire mdout1_5_13;
    wire mdout1_4_13;
    wire mdout1_3_13;
    wire mdout1_2_13;
    wire mdout1_1_13;
    wire mdout1_0_13;
    wire mdout1_7_14;
    wire mdout1_6_14;
    wire mdout1_5_14;
    wire mdout1_4_14;
    wire mdout1_3_14;
    wire mdout1_2_14;
    wire mdout1_1_14;
    wire mdout1_0_14;
    wire mdout1_7_15;
    wire mdout1_6_15;
    wire mdout1_5_15;
    wire mdout1_4_15;
    wire mdout1_3_15;
    wire mdout1_2_15;
    wire mdout1_1_15;
    wire mdout1_0_15;
    wire mdout1_7_16;
    wire mdout1_6_16;
    wire mdout1_5_16;
    wire mdout1_4_16;
    wire mdout1_3_16;
    wire mdout1_2_16;
    wire mdout1_1_16;
    wire mdout1_0_16;
    wire mdout1_7_17;
    wire mdout1_6_17;
    wire mdout1_5_17;
    wire mdout1_4_17;
    wire mdout1_3_17;
    wire mdout1_2_17;
    wire mdout1_1_17;
    wire mdout1_0_17;
    wire mdout1_7_18;
    wire mdout1_6_18;
    wire mdout1_5_18;
    wire mdout1_4_18;
    wire mdout1_3_18;
    wire mdout1_2_18;
    wire mdout1_1_18;
    wire mdout1_0_18;
    wire mdout1_7_19;
    wire mdout1_6_19;
    wire mdout1_5_19;
    wire mdout1_4_19;
    wire mdout1_3_19;
    wire mdout1_2_19;
    wire mdout1_1_19;
    wire mdout1_0_19;
    wire mdout1_7_20;
    wire mdout1_6_20;
    wire mdout1_5_20;
    wire mdout1_4_20;
    wire mdout1_3_20;
    wire mdout1_2_20;
    wire mdout1_1_20;
    wire mdout1_0_20;
    wire mdout1_7_21;
    wire mdout1_6_21;
    wire mdout1_5_21;
    wire mdout1_4_21;
    wire mdout1_3_21;
    wire mdout1_2_21;
    wire mdout1_1_21;
    wire mdout1_0_21;
    wire mdout1_7_22;
    wire mdout1_6_22;
    wire mdout1_5_22;
    wire mdout1_4_22;
    wire mdout1_3_22;
    wire mdout1_2_22;
    wire mdout1_1_22;
    wire mdout1_0_22;
    wire mdout1_7_23;
    wire mdout1_6_23;
    wire mdout1_5_23;
    wire mdout1_4_23;
    wire mdout1_3_23;
    wire mdout1_2_23;
    wire mdout1_1_23;
    wire mdout1_0_23;
    wire mdout1_7_24;
    wire mdout1_6_24;
    wire mdout1_5_24;
    wire mdout1_4_24;
    wire mdout1_3_24;
    wire mdout1_2_24;
    wire mdout1_1_24;
    wire mdout1_0_24;
    wire mdout1_7_25;
    wire mdout1_6_25;
    wire mdout1_5_25;
    wire mdout1_4_25;
    wire mdout1_3_25;
    wire mdout1_2_25;
    wire mdout1_1_25;
    wire mdout1_0_25;
    wire mdout1_7_26;
    wire mdout1_6_26;
    wire mdout1_5_26;
    wire mdout1_4_26;
    wire mdout1_3_26;
    wire mdout1_2_26;
    wire mdout1_1_26;
    wire mdout1_0_26;
    wire mdout1_7_27;
    wire mdout1_6_27;
    wire mdout1_5_27;
    wire mdout1_4_27;
    wire mdout1_3_27;
    wire mdout1_2_27;
    wire mdout1_1_27;
    wire mdout1_0_27;
    wire mdout1_7_28;
    wire mdout1_6_28;
    wire mdout1_5_28;
    wire mdout1_4_28;
    wire mdout1_3_28;
    wire mdout1_2_28;
    wire mdout1_1_28;
    wire mdout1_0_28;
    wire mdout1_7_29;
    wire mdout1_6_29;
    wire mdout1_5_29;
    wire mdout1_4_29;
    wire mdout1_3_29;
    wire mdout1_2_29;
    wire mdout1_1_29;
    wire mdout1_0_29;
    wire mdout1_7_30;
    wire mdout1_6_30;
    wire mdout1_5_30;
    wire mdout1_4_30;
    wire mdout1_3_30;
    wire mdout1_2_30;
    wire mdout1_1_30;
    wire mdout1_0_30;
    wire mdout1_7_31;
    wire mdout1_6_31;
    wire mdout1_5_31;
    wire mdout1_4_31;
    wire mdout1_3_31;
    wire mdout1_2_31;
    wire mdout1_1_31;
    wire mdout1_0_31;
    wire mdout1_7_32;
    wire mdout1_6_32;
    wire mdout1_5_32;
    wire mdout1_4_32;
    wire mdout1_3_32;
    wire mdout1_2_32;
    wire mdout1_1_32;
    wire mdout1_0_32;
    wire mdout1_7_33;
    wire mdout1_6_33;
    wire mdout1_5_33;
    wire mdout1_4_33;
    wire mdout1_3_33;
    wire mdout1_2_33;
    wire mdout1_1_33;
    wire mdout1_0_33;
    wire mdout1_7_34;
    wire mdout1_6_34;
    wire mdout1_5_34;
    wire mdout1_4_34;
    wire mdout1_3_34;
    wire mdout1_2_34;
    wire mdout1_1_34;
    wire mdout1_0_34;
    wire mdout1_7_35;
    wire mdout1_6_35;
    wire mdout1_5_35;
    wire mdout1_4_35;
    wire mdout1_3_35;
    wire mdout1_2_35;
    wire mdout1_1_35;
    wire mdout1_0_35;
    wire mdout1_7_36;
    wire mdout1_6_36;
    wire mdout1_5_36;
    wire mdout1_4_36;
    wire mdout1_3_36;
    wire mdout1_2_36;
    wire mdout1_1_36;
    wire mdout1_0_36;
    wire mdout1_7_37;
    wire mdout1_6_37;
    wire mdout1_5_37;
    wire mdout1_4_37;
    wire mdout1_3_37;
    wire mdout1_2_37;
    wire mdout1_1_37;
    wire mdout1_0_37;
    wire mdout1_7_38;
    wire mdout1_6_38;
    wire mdout1_5_38;
    wire mdout1_4_38;
    wire mdout1_3_38;
    wire mdout1_2_38;
    wire mdout1_1_38;
    wire mdout1_0_38;
    wire mdout1_7_39;
    wire mdout1_6_39;
    wire mdout1_5_39;
    wire mdout1_4_39;
    wire mdout1_3_39;
    wire mdout1_2_39;
    wire mdout1_1_39;
    wire mdout1_0_39;
    wire mdout1_7_40;
    wire mdout1_6_40;
    wire mdout1_5_40;
    wire mdout1_4_40;
    wire mdout1_3_40;
    wire mdout1_2_40;
    wire mdout1_1_40;
    wire mdout1_0_40;
    wire mdout1_7_41;
    wire mdout1_6_41;
    wire mdout1_5_41;
    wire mdout1_4_41;
    wire mdout1_3_41;
    wire mdout1_2_41;
    wire mdout1_1_41;
    wire mdout1_0_41;
    wire mdout1_7_42;
    wire mdout1_6_42;
    wire mdout1_5_42;
    wire mdout1_4_42;
    wire mdout1_3_42;
    wire mdout1_2_42;
    wire mdout1_1_42;
    wire mdout1_0_42;
    wire mdout1_7_43;
    wire mdout1_6_43;
    wire mdout1_5_43;
    wire mdout1_4_43;
    wire mdout1_3_43;
    wire mdout1_2_43;
    wire mdout1_1_43;
    wire mdout1_0_43;
    wire mdout1_7_44;
    wire mdout1_6_44;
    wire mdout1_5_44;
    wire mdout1_4_44;
    wire mdout1_3_44;
    wire mdout1_2_44;
    wire mdout1_1_44;
    wire mdout1_0_44;
    wire mdout1_7_45;
    wire mdout1_6_45;
    wire mdout1_5_45;
    wire mdout1_4_45;
    wire mdout1_3_45;
    wire mdout1_2_45;
    wire mdout1_1_45;
    wire mdout1_0_45;
    wire mdout1_7_46;
    wire mdout1_6_46;
    wire mdout1_5_46;
    wire mdout1_4_46;
    wire mdout1_3_46;
    wire mdout1_2_46;
    wire mdout1_1_46;
    wire mdout1_0_46;
    wire mdout1_7_47;
    wire mdout1_6_47;
    wire mdout1_5_47;
    wire mdout1_4_47;
    wire mdout1_3_47;
    wire mdout1_2_47;
    wire mdout1_1_47;
    wire mdout1_0_47;
    wire mdout1_7_48;
    wire mdout1_6_48;
    wire mdout1_5_48;
    wire mdout1_4_48;
    wire mdout1_3_48;
    wire mdout1_2_48;
    wire mdout1_1_48;
    wire mdout1_0_48;
    wire mdout1_7_49;
    wire mdout1_6_49;
    wire mdout1_5_49;
    wire mdout1_4_49;
    wire mdout1_3_49;
    wire mdout1_2_49;
    wire mdout1_1_49;
    wire mdout1_0_49;
    wire mdout1_7_50;
    wire mdout1_6_50;
    wire mdout1_5_50;
    wire mdout1_4_50;
    wire mdout1_3_50;
    wire mdout1_2_50;
    wire mdout1_1_50;
    wire mdout1_0_50;
    wire mdout1_7_51;
    wire mdout1_6_51;
    wire mdout1_5_51;
    wire mdout1_4_51;
    wire mdout1_3_51;
    wire mdout1_2_51;
    wire mdout1_1_51;
    wire mdout1_0_51;
    wire mdout1_7_52;
    wire mdout1_6_52;
    wire mdout1_5_52;
    wire mdout1_4_52;
    wire mdout1_3_52;
    wire mdout1_2_52;
    wire mdout1_1_52;
    wire mdout1_0_52;
    wire mdout1_7_53;
    wire mdout1_6_53;
    wire mdout1_5_53;
    wire mdout1_4_53;
    wire mdout1_3_53;
    wire mdout1_2_53;
    wire mdout1_1_53;
    wire mdout1_0_53;
    wire mdout1_7_54;
    wire mdout1_6_54;
    wire mdout1_5_54;
    wire mdout1_4_54;
    wire mdout1_3_54;
    wire mdout1_2_54;
    wire mdout1_1_54;
    wire mdout1_0_54;
    wire mdout1_7_55;
    wire mdout1_6_55;
    wire mdout1_5_55;
    wire mdout1_4_55;
    wire mdout1_3_55;
    wire mdout1_2_55;
    wire mdout1_1_55;
    wire mdout1_0_55;
    wire mdout1_7_56;
    wire mdout1_6_56;
    wire mdout1_5_56;
    wire mdout1_4_56;
    wire mdout1_3_56;
    wire mdout1_2_56;
    wire mdout1_1_56;
    wire mdout1_0_56;
    wire mdout1_7_57;
    wire mdout1_6_57;
    wire mdout1_5_57;
    wire mdout1_4_57;
    wire mdout1_3_57;
    wire mdout1_2_57;
    wire mdout1_1_57;
    wire mdout1_0_57;
    wire mdout1_7_58;
    wire mdout1_6_58;
    wire mdout1_5_58;
    wire mdout1_4_58;
    wire mdout1_3_58;
    wire mdout1_2_58;
    wire mdout1_1_58;
    wire mdout1_0_58;
    wire mdout1_7_59;
    wire mdout1_6_59;
    wire mdout1_5_59;
    wire mdout1_4_59;
    wire mdout1_3_59;
    wire mdout1_2_59;
    wire mdout1_1_59;
    wire mdout1_0_59;
    wire mdout1_7_60;
    wire mdout1_6_60;
    wire mdout1_5_60;
    wire mdout1_4_60;
    wire mdout1_3_60;
    wire mdout1_2_60;
    wire mdout1_1_60;
    wire mdout1_0_60;
    wire mdout1_7_61;
    wire mdout1_6_61;
    wire mdout1_5_61;
    wire mdout1_4_61;
    wire mdout1_3_61;
    wire mdout1_2_61;
    wire mdout1_1_61;
    wire mdout1_0_61;
    wire mdout1_7_62;
    wire mdout1_6_62;
    wire mdout1_5_62;
    wire mdout1_4_62;
    wire mdout1_3_62;
    wire mdout1_2_62;
    wire mdout1_1_62;
    wire mdout1_0_62;
    wire mdout1_7_63;
    wire mdout1_6_63;
    wire mdout1_5_63;
    wire mdout1_4_63;
    wire mdout1_3_63;
    wire mdout1_2_63;
    wire mdout1_1_63;
    wire mdout1_0_63;
    wire mdout1_7_64;
    wire mdout1_6_64;
    wire mdout1_5_64;
    wire mdout1_4_64;
    wire mdout1_3_64;
    wire mdout1_2_64;
    wire mdout1_1_64;
    wire mdout1_0_64;
    wire mdout1_7_65;
    wire mdout1_6_65;
    wire mdout1_5_65;
    wire mdout1_4_65;
    wire mdout1_3_65;
    wire mdout1_2_65;
    wire mdout1_1_65;
    wire mdout1_0_65;
    wire mdout1_7_66;
    wire mdout1_6_66;
    wire mdout1_5_66;
    wire mdout1_4_66;
    wire mdout1_3_66;
    wire mdout1_2_66;
    wire mdout1_1_66;
    wire mdout1_0_66;
    wire mdout1_7_67;
    wire mdout1_6_67;
    wire mdout1_5_67;
    wire mdout1_4_67;
    wire mdout1_3_67;
    wire mdout1_2_67;
    wire mdout1_1_67;
    wire mdout1_0_67;
    wire mdout1_7_68;
    wire mdout1_6_68;
    wire mdout1_5_68;
    wire mdout1_4_68;
    wire mdout1_3_68;
    wire mdout1_2_68;
    wire mdout1_1_68;
    wire mdout1_0_68;
    wire mdout1_7_69;
    wire mdout1_6_69;
    wire mdout1_5_69;
    wire mdout1_4_69;
    wire mdout1_3_69;
    wire mdout1_2_69;
    wire mdout1_1_69;
    wire mdout1_0_69;
    wire mdout1_7_70;
    wire mdout1_6_70;
    wire mdout1_5_70;
    wire mdout1_4_70;
    wire mdout1_3_70;
    wire mdout1_2_70;
    wire mdout1_1_70;
    wire mdout1_0_70;
    wire mdout1_7_71;
    wire mdout1_6_71;
    wire mdout1_5_71;
    wire mdout1_4_71;
    wire mdout1_3_71;
    wire mdout1_2_71;
    wire mdout1_1_71;
    wire mdout1_0_71;
    wire mdout1_7_72;
    wire mdout1_6_72;
    wire mdout1_5_72;
    wire mdout1_4_72;
    wire mdout1_3_72;
    wire mdout1_2_72;
    wire mdout1_1_72;
    wire mdout1_0_72;
    wire mdout1_7_73;
    wire mdout1_6_73;
    wire mdout1_5_73;
    wire mdout1_4_73;
    wire mdout1_3_73;
    wire mdout1_2_73;
    wire mdout1_1_73;
    wire mdout1_0_73;
    wire mdout1_7_74;
    wire mdout1_6_74;
    wire mdout1_5_74;
    wire mdout1_4_74;
    wire mdout1_3_74;
    wire mdout1_2_74;
    wire mdout1_1_74;
    wire mdout1_0_74;
    wire mdout1_7_75;
    wire mdout1_6_75;
    wire mdout1_5_75;
    wire mdout1_4_75;
    wire mdout1_3_75;
    wire mdout1_2_75;
    wire mdout1_1_75;
    wire mdout1_0_75;
    wire mdout1_7_76;
    wire mdout1_6_76;
    wire mdout1_5_76;
    wire mdout1_4_76;
    wire mdout1_3_76;
    wire mdout1_2_76;
    wire mdout1_1_76;
    wire mdout1_0_76;
    wire mdout1_7_77;
    wire mdout1_6_77;
    wire mdout1_5_77;
    wire mdout1_4_77;
    wire mdout1_3_77;
    wire mdout1_2_77;
    wire mdout1_1_77;
    wire mdout1_0_77;
    wire mdout1_7_78;
    wire mdout1_6_78;
    wire mdout1_5_78;
    wire mdout1_4_78;
    wire mdout1_3_78;
    wire mdout1_2_78;
    wire mdout1_1_78;
    wire mdout1_0_78;
    wire mdout1_7_79;
    wire mdout1_6_79;
    wire mdout1_5_79;
    wire mdout1_4_79;
    wire mdout1_3_79;
    wire mdout1_2_79;
    wire mdout1_1_79;
    wire mdout1_0_79;
    wire mdout1_7_80;
    wire mdout1_6_80;
    wire mdout1_5_80;
    wire mdout1_4_80;
    wire mdout1_3_80;
    wire mdout1_2_80;
    wire mdout1_1_80;
    wire mdout1_0_80;
    wire mdout1_7_81;
    wire mdout1_6_81;
    wire mdout1_5_81;
    wire mdout1_4_81;
    wire mdout1_3_81;
    wire mdout1_2_81;
    wire mdout1_1_81;
    wire mdout1_0_81;
    wire mdout1_7_82;
    wire mdout1_6_82;
    wire mdout1_5_82;
    wire mdout1_4_82;
    wire mdout1_3_82;
    wire mdout1_2_82;
    wire mdout1_1_82;
    wire mdout1_0_82;
    wire mdout1_7_83;
    wire mdout1_6_83;
    wire mdout1_5_83;
    wire mdout1_4_83;
    wire mdout1_3_83;
    wire mdout1_2_83;
    wire mdout1_1_83;
    wire mdout1_0_83;
    wire mdout1_7_84;
    wire mdout1_6_84;
    wire mdout1_5_84;
    wire mdout1_4_84;
    wire mdout1_3_84;
    wire mdout1_2_84;
    wire mdout1_1_84;
    wire mdout1_0_84;
    wire mdout1_7_85;
    wire mdout1_6_85;
    wire mdout1_5_85;
    wire mdout1_4_85;
    wire mdout1_3_85;
    wire mdout1_2_85;
    wire mdout1_1_85;
    wire mdout1_0_85;
    wire mdout1_7_86;
    wire mdout1_6_86;
    wire mdout1_5_86;
    wire mdout1_4_86;
    wire mdout1_3_86;
    wire mdout1_2_86;
    wire mdout1_1_86;
    wire mdout1_0_86;
    wire mdout1_7_87;
    wire mdout1_6_87;
    wire mdout1_5_87;
    wire mdout1_4_87;
    wire mdout1_3_87;
    wire mdout1_2_87;
    wire mdout1_1_87;
    wire mdout1_0_87;
    wire mdout1_7_88;
    wire mdout1_6_88;
    wire mdout1_5_88;
    wire mdout1_4_88;
    wire mdout1_3_88;
    wire mdout1_2_88;
    wire mdout1_1_88;
    wire mdout1_0_88;
    wire mdout1_7_89;
    wire mdout1_6_89;
    wire mdout1_5_89;
    wire mdout1_4_89;
    wire mdout1_3_89;
    wire mdout1_2_89;
    wire mdout1_1_89;
    wire mdout1_0_89;
    wire mdout1_7_90;
    wire mdout1_6_90;
    wire mdout1_5_90;
    wire mdout1_4_90;
    wire mdout1_3_90;
    wire mdout1_2_90;
    wire mdout1_1_90;
    wire mdout1_0_90;
    wire mdout1_7_91;
    wire mdout1_6_91;
    wire mdout1_5_91;
    wire mdout1_4_91;
    wire mdout1_3_91;
    wire mdout1_2_91;
    wire mdout1_1_91;
    wire mdout1_0_91;
    wire mdout1_7_92;
    wire mdout1_6_92;
    wire mdout1_5_92;
    wire mdout1_4_92;
    wire mdout1_3_92;
    wire mdout1_2_92;
    wire mdout1_1_92;
    wire mdout1_0_92;
    wire mdout1_7_93;
    wire mdout1_6_93;
    wire mdout1_5_93;
    wire mdout1_4_93;
    wire mdout1_3_93;
    wire mdout1_2_93;
    wire mdout1_1_93;
    wire mdout1_0_93;
    wire mdout1_7_94;
    wire mdout1_6_94;
    wire mdout1_5_94;
    wire mdout1_4_94;
    wire mdout1_3_94;
    wire mdout1_2_94;
    wire mdout1_1_94;
    wire mdout1_0_94;
    wire mdout1_7_95;
    wire mdout1_6_95;
    wire mdout1_5_95;
    wire mdout1_4_95;
    wire mdout1_3_95;
    wire mdout1_2_95;
    wire mdout1_1_95;
    wire mdout1_0_95;
    wire mdout1_7_96;
    wire mdout1_6_96;
    wire mdout1_5_96;
    wire mdout1_4_96;
    wire mdout1_3_96;
    wire mdout1_2_96;
    wire mdout1_1_96;
    wire mdout1_0_96;
    wire mdout1_7_97;
    wire mdout1_6_97;
    wire mdout1_5_97;
    wire mdout1_4_97;
    wire mdout1_3_97;
    wire mdout1_2_97;
    wire mdout1_1_97;
    wire mdout1_0_97;
    wire raddr13_ff2;
    wire raddr12_ff2;
    wire raddr11_ff2;
    wire mdout1_7_98;
    wire mdout1_6_98;
    wire mdout1_5_98;
    wire mdout1_4_98;
    wire mdout1_3_98;
    wire mdout1_2_98;
    wire mdout1_1_98;
    wire mdout1_0_98;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87 (.DIA0(Data[0]), 
        .DIA1(Data[1]), .DIA2(Data[2]), .DIA3(Data[3]), .DIA4(Data[4]), 
        .DIA5(Data[5]), .DIA6(Data[6]), .DIA7(Data[7]), .DIA8(Data[8]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_0), 
        .DOB1(mdout1_0_1), .DOB2(mdout1_0_2), .DOB3(mdout1_0_3), .DOB4(mdout1_0_4), 
        .DOB5(mdout1_0_5), .DOB6(mdout1_0_6), .DOB7(mdout1_0_7), .DOB8(mdout1_0_8), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86 (.DIA0(Data[9]), 
        .DIA1(Data[10]), .DIA2(Data[11]), .DIA3(Data[12]), .DIA4(Data[13]), 
        .DIA5(Data[14]), .DIA6(Data[15]), .DIA7(Data[16]), .DIA8(Data[17]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_9), 
        .DOB1(mdout1_0_10), .DOB2(mdout1_0_11), .DOB3(mdout1_0_12), .DOB4(mdout1_0_13), 
        .DOB5(mdout1_0_14), .DOB6(mdout1_0_15), .DOB7(mdout1_0_16), .DOB8(mdout1_0_17), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85 (.DIA0(Data[18]), 
        .DIA1(Data[19]), .DIA2(Data[20]), .DIA3(Data[21]), .DIA4(Data[22]), 
        .DIA5(Data[23]), .DIA6(Data[24]), .DIA7(Data[25]), .DIA8(Data[26]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_18), 
        .DOB1(mdout1_0_19), .DOB2(mdout1_0_20), .DOB3(mdout1_0_21), .DOB4(mdout1_0_22), 
        .DOB5(mdout1_0_23), .DOB6(mdout1_0_24), .DOB7(mdout1_0_25), .DOB8(mdout1_0_26), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84 (.DIA0(Data[27]), 
        .DIA1(Data[28]), .DIA2(Data[29]), .DIA3(Data[30]), .DIA4(Data[31]), 
        .DIA5(Data[32]), .DIA6(Data[33]), .DIA7(Data[34]), .DIA8(Data[35]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_27), 
        .DOB1(mdout1_0_28), .DOB2(mdout1_0_29), .DOB3(mdout1_0_30), .DOB4(mdout1_0_31), 
        .DOB5(mdout1_0_32), .DOB6(mdout1_0_33), .DOB7(mdout1_0_34), .DOB8(mdout1_0_35), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83 (.DIA0(Data[36]), 
        .DIA1(Data[37]), .DIA2(Data[38]), .DIA3(Data[39]), .DIA4(Data[40]), 
        .DIA5(Data[41]), .DIA6(Data[42]), .DIA7(Data[43]), .DIA8(Data[44]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_36), 
        .DOB1(mdout1_0_37), .DOB2(mdout1_0_38), .DOB3(mdout1_0_39), .DOB4(mdout1_0_40), 
        .DOB5(mdout1_0_41), .DOB6(mdout1_0_42), .DOB7(mdout1_0_43), .DOB8(mdout1_0_44), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82 (.DIA0(Data[45]), 
        .DIA1(Data[46]), .DIA2(Data[47]), .DIA3(Data[48]), .DIA4(Data[49]), 
        .DIA5(Data[50]), .DIA6(Data[51]), .DIA7(Data[52]), .DIA8(Data[53]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_45), 
        .DOB1(mdout1_0_46), .DOB2(mdout1_0_47), .DOB3(mdout1_0_48), .DOB4(mdout1_0_49), 
        .DOB5(mdout1_0_50), .DOB6(mdout1_0_51), .DOB7(mdout1_0_52), .DOB8(mdout1_0_53), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81 (.DIA0(Data[54]), 
        .DIA1(Data[55]), .DIA2(Data[56]), .DIA3(Data[57]), .DIA4(Data[58]), 
        .DIA5(Data[59]), .DIA6(Data[60]), .DIA7(Data[61]), .DIA8(Data[62]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_54), 
        .DOB1(mdout1_0_55), .DOB2(mdout1_0_56), .DOB3(mdout1_0_57), .DOB4(mdout1_0_58), 
        .DOB5(mdout1_0_59), .DOB6(mdout1_0_60), .DOB7(mdout1_0_61), .DOB8(mdout1_0_62), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80 (.DIA0(Data[63]), 
        .DIA1(Data[64]), .DIA2(Data[65]), .DIA3(Data[66]), .DIA4(Data[67]), 
        .DIA5(Data[68]), .DIA6(Data[69]), .DIA7(Data[70]), .DIA8(Data[71]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_63), 
        .DOB1(mdout1_0_64), .DOB2(mdout1_0_65), .DOB3(mdout1_0_66), .DOB4(mdout1_0_67), 
        .DOB5(mdout1_0_68), .DOB6(mdout1_0_69), .DOB7(mdout1_0_70), .DOB8(mdout1_0_71), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79 (.DIA0(Data[72]), 
        .DIA1(Data[73]), .DIA2(Data[74]), .DIA3(Data[75]), .DIA4(Data[76]), 
        .DIA5(Data[77]), .DIA6(Data[78]), .DIA7(Data[79]), .DIA8(Data[80]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_72), 
        .DOB1(mdout1_0_73), .DOB2(mdout1_0_74), .DOB3(mdout1_0_75), .DOB4(mdout1_0_76), 
        .DOB5(mdout1_0_77), .DOB6(mdout1_0_78), .DOB7(mdout1_0_79), .DOB8(mdout1_0_80), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78 (.DIA0(Data[81]), 
        .DIA1(Data[82]), .DIA2(Data[83]), .DIA3(Data[84]), .DIA4(Data[85]), 
        .DIA5(Data[86]), .DIA6(Data[87]), .DIA7(Data[88]), .DIA8(Data[89]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_81), 
        .DOB1(mdout1_0_82), .DOB2(mdout1_0_83), .DOB3(mdout1_0_84), .DOB4(mdout1_0_85), 
        .DOB5(mdout1_0_86), .DOB6(mdout1_0_87), .DOB7(mdout1_0_88), .DOB8(mdout1_0_89), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77 (.DIA0(Data[90]), 
        .DIA1(Data[91]), .DIA2(Data[92]), .DIA3(Data[93]), .DIA4(Data[94]), 
        .DIA5(Data[95]), .DIA6(Data[96]), .DIA7(Data[97]), .DIA8(Data[98]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_0_90), 
        .DOB1(mdout1_0_91), .DOB2(mdout1_0_92), .DOB3(mdout1_0_93), .DOB4(mdout1_0_94), 
        .DOB5(mdout1_0_95), .DOB6(mdout1_0_96), .DOB7(mdout1_0_97), .DOB8(mdout1_0_98), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76 (.DIA0(Data[0]), 
        .DIA1(Data[1]), .DIA2(Data[2]), .DIA3(Data[3]), .DIA4(Data[4]), 
        .DIA5(Data[5]), .DIA6(Data[6]), .DIA7(Data[7]), .DIA8(Data[8]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_0), 
        .DOB1(mdout1_1_1), .DOB2(mdout1_1_2), .DOB3(mdout1_1_3), .DOB4(mdout1_1_4), 
        .DOB5(mdout1_1_5), .DOB6(mdout1_1_6), .DOB7(mdout1_1_7), .DOB8(mdout1_1_8), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75 (.DIA0(Data[9]), 
        .DIA1(Data[10]), .DIA2(Data[11]), .DIA3(Data[12]), .DIA4(Data[13]), 
        .DIA5(Data[14]), .DIA6(Data[15]), .DIA7(Data[16]), .DIA8(Data[17]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_9), 
        .DOB1(mdout1_1_10), .DOB2(mdout1_1_11), .DOB3(mdout1_1_12), .DOB4(mdout1_1_13), 
        .DOB5(mdout1_1_14), .DOB6(mdout1_1_15), .DOB7(mdout1_1_16), .DOB8(mdout1_1_17), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74 (.DIA0(Data[18]), 
        .DIA1(Data[19]), .DIA2(Data[20]), .DIA3(Data[21]), .DIA4(Data[22]), 
        .DIA5(Data[23]), .DIA6(Data[24]), .DIA7(Data[25]), .DIA8(Data[26]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_18), 
        .DOB1(mdout1_1_19), .DOB2(mdout1_1_20), .DOB3(mdout1_1_21), .DOB4(mdout1_1_22), 
        .DOB5(mdout1_1_23), .DOB6(mdout1_1_24), .DOB7(mdout1_1_25), .DOB8(mdout1_1_26), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73 (.DIA0(Data[27]), 
        .DIA1(Data[28]), .DIA2(Data[29]), .DIA3(Data[30]), .DIA4(Data[31]), 
        .DIA5(Data[32]), .DIA6(Data[33]), .DIA7(Data[34]), .DIA8(Data[35]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_27), 
        .DOB1(mdout1_1_28), .DOB2(mdout1_1_29), .DOB3(mdout1_1_30), .DOB4(mdout1_1_31), 
        .DOB5(mdout1_1_32), .DOB6(mdout1_1_33), .DOB7(mdout1_1_34), .DOB8(mdout1_1_35), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72 (.DIA0(Data[36]), 
        .DIA1(Data[37]), .DIA2(Data[38]), .DIA3(Data[39]), .DIA4(Data[40]), 
        .DIA5(Data[41]), .DIA6(Data[42]), .DIA7(Data[43]), .DIA8(Data[44]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_36), 
        .DOB1(mdout1_1_37), .DOB2(mdout1_1_38), .DOB3(mdout1_1_39), .DOB4(mdout1_1_40), 
        .DOB5(mdout1_1_41), .DOB6(mdout1_1_42), .DOB7(mdout1_1_43), .DOB8(mdout1_1_44), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71 (.DIA0(Data[45]), 
        .DIA1(Data[46]), .DIA2(Data[47]), .DIA3(Data[48]), .DIA4(Data[49]), 
        .DIA5(Data[50]), .DIA6(Data[51]), .DIA7(Data[52]), .DIA8(Data[53]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_45), 
        .DOB1(mdout1_1_46), .DOB2(mdout1_1_47), .DOB3(mdout1_1_48), .DOB4(mdout1_1_49), 
        .DOB5(mdout1_1_50), .DOB6(mdout1_1_51), .DOB7(mdout1_1_52), .DOB8(mdout1_1_53), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70 (.DIA0(Data[54]), 
        .DIA1(Data[55]), .DIA2(Data[56]), .DIA3(Data[57]), .DIA4(Data[58]), 
        .DIA5(Data[59]), .DIA6(Data[60]), .DIA7(Data[61]), .DIA8(Data[62]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_54), 
        .DOB1(mdout1_1_55), .DOB2(mdout1_1_56), .DOB3(mdout1_1_57), .DOB4(mdout1_1_58), 
        .DOB5(mdout1_1_59), .DOB6(mdout1_1_60), .DOB7(mdout1_1_61), .DOB8(mdout1_1_62), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69 (.DIA0(Data[63]), 
        .DIA1(Data[64]), .DIA2(Data[65]), .DIA3(Data[66]), .DIA4(Data[67]), 
        .DIA5(Data[68]), .DIA6(Data[69]), .DIA7(Data[70]), .DIA8(Data[71]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_63), 
        .DOB1(mdout1_1_64), .DOB2(mdout1_1_65), .DOB3(mdout1_1_66), .DOB4(mdout1_1_67), 
        .DOB5(mdout1_1_68), .DOB6(mdout1_1_69), .DOB7(mdout1_1_70), .DOB8(mdout1_1_71), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68 (.DIA0(Data[72]), 
        .DIA1(Data[73]), .DIA2(Data[74]), .DIA3(Data[75]), .DIA4(Data[76]), 
        .DIA5(Data[77]), .DIA6(Data[78]), .DIA7(Data[79]), .DIA8(Data[80]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_72), 
        .DOB1(mdout1_1_73), .DOB2(mdout1_1_74), .DOB3(mdout1_1_75), .DOB4(mdout1_1_76), 
        .DOB5(mdout1_1_77), .DOB6(mdout1_1_78), .DOB7(mdout1_1_79), .DOB8(mdout1_1_80), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67 (.DIA0(Data[81]), 
        .DIA1(Data[82]), .DIA2(Data[83]), .DIA3(Data[84]), .DIA4(Data[85]), 
        .DIA5(Data[86]), .DIA6(Data[87]), .DIA7(Data[88]), .DIA8(Data[89]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_81), 
        .DOB1(mdout1_1_82), .DOB2(mdout1_1_83), .DOB3(mdout1_1_84), .DOB4(mdout1_1_85), 
        .DOB5(mdout1_1_86), .DOB6(mdout1_1_87), .DOB7(mdout1_1_88), .DOB8(mdout1_1_89), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66 (.DIA0(Data[90]), 
        .DIA1(Data[91]), .DIA2(Data[92]), .DIA3(Data[93]), .DIA4(Data[94]), 
        .DIA5(Data[95]), .DIA6(Data[96]), .DIA7(Data[97]), .DIA8(Data[98]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_1_90), 
        .DOB1(mdout1_1_91), .DOB2(mdout1_1_92), .DOB3(mdout1_1_93), .DOB4(mdout1_1_94), 
        .DOB5(mdout1_1_95), .DOB6(mdout1_1_96), .DOB7(mdout1_1_97), .DOB8(mdout1_1_98), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65 (.DIA0(Data[0]), 
        .DIA1(Data[1]), .DIA2(Data[2]), .DIA3(Data[3]), .DIA4(Data[4]), 
        .DIA5(Data[5]), .DIA6(Data[6]), .DIA7(Data[7]), .DIA8(Data[8]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_0), 
        .DOB1(mdout1_2_1), .DOB2(mdout1_2_2), .DOB3(mdout1_2_3), .DOB4(mdout1_2_4), 
        .DOB5(mdout1_2_5), .DOB6(mdout1_2_6), .DOB7(mdout1_2_7), .DOB8(mdout1_2_8), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64 (.DIA0(Data[9]), 
        .DIA1(Data[10]), .DIA2(Data[11]), .DIA3(Data[12]), .DIA4(Data[13]), 
        .DIA5(Data[14]), .DIA6(Data[15]), .DIA7(Data[16]), .DIA8(Data[17]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_9), 
        .DOB1(mdout1_2_10), .DOB2(mdout1_2_11), .DOB3(mdout1_2_12), .DOB4(mdout1_2_13), 
        .DOB5(mdout1_2_14), .DOB6(mdout1_2_15), .DOB7(mdout1_2_16), .DOB8(mdout1_2_17), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63 (.DIA0(Data[18]), 
        .DIA1(Data[19]), .DIA2(Data[20]), .DIA3(Data[21]), .DIA4(Data[22]), 
        .DIA5(Data[23]), .DIA6(Data[24]), .DIA7(Data[25]), .DIA8(Data[26]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_18), 
        .DOB1(mdout1_2_19), .DOB2(mdout1_2_20), .DOB3(mdout1_2_21), .DOB4(mdout1_2_22), 
        .DOB5(mdout1_2_23), .DOB6(mdout1_2_24), .DOB7(mdout1_2_25), .DOB8(mdout1_2_26), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62 (.DIA0(Data[27]), 
        .DIA1(Data[28]), .DIA2(Data[29]), .DIA3(Data[30]), .DIA4(Data[31]), 
        .DIA5(Data[32]), .DIA6(Data[33]), .DIA7(Data[34]), .DIA8(Data[35]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_27), 
        .DOB1(mdout1_2_28), .DOB2(mdout1_2_29), .DOB3(mdout1_2_30), .DOB4(mdout1_2_31), 
        .DOB5(mdout1_2_32), .DOB6(mdout1_2_33), .DOB7(mdout1_2_34), .DOB8(mdout1_2_35), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61 (.DIA0(Data[36]), 
        .DIA1(Data[37]), .DIA2(Data[38]), .DIA3(Data[39]), .DIA4(Data[40]), 
        .DIA5(Data[41]), .DIA6(Data[42]), .DIA7(Data[43]), .DIA8(Data[44]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_36), 
        .DOB1(mdout1_2_37), .DOB2(mdout1_2_38), .DOB3(mdout1_2_39), .DOB4(mdout1_2_40), 
        .DOB5(mdout1_2_41), .DOB6(mdout1_2_42), .DOB7(mdout1_2_43), .DOB8(mdout1_2_44), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60 (.DIA0(Data[45]), 
        .DIA1(Data[46]), .DIA2(Data[47]), .DIA3(Data[48]), .DIA4(Data[49]), 
        .DIA5(Data[50]), .DIA6(Data[51]), .DIA7(Data[52]), .DIA8(Data[53]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_45), 
        .DOB1(mdout1_2_46), .DOB2(mdout1_2_47), .DOB3(mdout1_2_48), .DOB4(mdout1_2_49), 
        .DOB5(mdout1_2_50), .DOB6(mdout1_2_51), .DOB7(mdout1_2_52), .DOB8(mdout1_2_53), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59 (.DIA0(Data[54]), 
        .DIA1(Data[55]), .DIA2(Data[56]), .DIA3(Data[57]), .DIA4(Data[58]), 
        .DIA5(Data[59]), .DIA6(Data[60]), .DIA7(Data[61]), .DIA8(Data[62]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_54), 
        .DOB1(mdout1_2_55), .DOB2(mdout1_2_56), .DOB3(mdout1_2_57), .DOB4(mdout1_2_58), 
        .DOB5(mdout1_2_59), .DOB6(mdout1_2_60), .DOB7(mdout1_2_61), .DOB8(mdout1_2_62), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58 (.DIA0(Data[63]), 
        .DIA1(Data[64]), .DIA2(Data[65]), .DIA3(Data[66]), .DIA4(Data[67]), 
        .DIA5(Data[68]), .DIA6(Data[69]), .DIA7(Data[70]), .DIA8(Data[71]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_63), 
        .DOB1(mdout1_2_64), .DOB2(mdout1_2_65), .DOB3(mdout1_2_66), .DOB4(mdout1_2_67), 
        .DOB5(mdout1_2_68), .DOB6(mdout1_2_69), .DOB7(mdout1_2_70), .DOB8(mdout1_2_71), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57 (.DIA0(Data[72]), 
        .DIA1(Data[73]), .DIA2(Data[74]), .DIA3(Data[75]), .DIA4(Data[76]), 
        .DIA5(Data[77]), .DIA6(Data[78]), .DIA7(Data[79]), .DIA8(Data[80]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_72), 
        .DOB1(mdout1_2_73), .DOB2(mdout1_2_74), .DOB3(mdout1_2_75), .DOB4(mdout1_2_76), 
        .DOB5(mdout1_2_77), .DOB6(mdout1_2_78), .DOB7(mdout1_2_79), .DOB8(mdout1_2_80), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56 (.DIA0(Data[81]), 
        .DIA1(Data[82]), .DIA2(Data[83]), .DIA3(Data[84]), .DIA4(Data[85]), 
        .DIA5(Data[86]), .DIA6(Data[87]), .DIA7(Data[88]), .DIA8(Data[89]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_81), 
        .DOB1(mdout1_2_82), .DOB2(mdout1_2_83), .DOB3(mdout1_2_84), .DOB4(mdout1_2_85), 
        .DOB5(mdout1_2_86), .DOB6(mdout1_2_87), .DOB7(mdout1_2_88), .DOB8(mdout1_2_89), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55.CSDECODE_B = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55.CSDECODE_A = "0b010" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55 (.DIA0(Data[90]), 
        .DIA1(Data[91]), .DIA2(Data[92]), .DIA3(Data[93]), .DIA4(Data[94]), 
        .DIA5(Data[95]), .DIA6(Data[96]), .DIA7(Data[97]), .DIA8(Data[98]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_2_90), 
        .DOB1(mdout1_2_91), .DOB2(mdout1_2_92), .DOB3(mdout1_2_93), .DOB4(mdout1_2_94), 
        .DOB5(mdout1_2_95), .DOB6(mdout1_2_96), .DOB7(mdout1_2_97), .DOB8(mdout1_2_98), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54 (.DIA0(Data[0]), 
        .DIA1(Data[1]), .DIA2(Data[2]), .DIA3(Data[3]), .DIA4(Data[4]), 
        .DIA5(Data[5]), .DIA6(Data[6]), .DIA7(Data[7]), .DIA8(Data[8]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_0), 
        .DOB1(mdout1_3_1), .DOB2(mdout1_3_2), .DOB3(mdout1_3_3), .DOB4(mdout1_3_4), 
        .DOB5(mdout1_3_5), .DOB6(mdout1_3_6), .DOB7(mdout1_3_7), .DOB8(mdout1_3_8), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53 (.DIA0(Data[9]), 
        .DIA1(Data[10]), .DIA2(Data[11]), .DIA3(Data[12]), .DIA4(Data[13]), 
        .DIA5(Data[14]), .DIA6(Data[15]), .DIA7(Data[16]), .DIA8(Data[17]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_9), 
        .DOB1(mdout1_3_10), .DOB2(mdout1_3_11), .DOB3(mdout1_3_12), .DOB4(mdout1_3_13), 
        .DOB5(mdout1_3_14), .DOB6(mdout1_3_15), .DOB7(mdout1_3_16), .DOB8(mdout1_3_17), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52 (.DIA0(Data[18]), 
        .DIA1(Data[19]), .DIA2(Data[20]), .DIA3(Data[21]), .DIA4(Data[22]), 
        .DIA5(Data[23]), .DIA6(Data[24]), .DIA7(Data[25]), .DIA8(Data[26]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_18), 
        .DOB1(mdout1_3_19), .DOB2(mdout1_3_20), .DOB3(mdout1_3_21), .DOB4(mdout1_3_22), 
        .DOB5(mdout1_3_23), .DOB6(mdout1_3_24), .DOB7(mdout1_3_25), .DOB8(mdout1_3_26), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51 (.DIA0(Data[27]), 
        .DIA1(Data[28]), .DIA2(Data[29]), .DIA3(Data[30]), .DIA4(Data[31]), 
        .DIA5(Data[32]), .DIA6(Data[33]), .DIA7(Data[34]), .DIA8(Data[35]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_27), 
        .DOB1(mdout1_3_28), .DOB2(mdout1_3_29), .DOB3(mdout1_3_30), .DOB4(mdout1_3_31), 
        .DOB5(mdout1_3_32), .DOB6(mdout1_3_33), .DOB7(mdout1_3_34), .DOB8(mdout1_3_35), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50 (.DIA0(Data[36]), 
        .DIA1(Data[37]), .DIA2(Data[38]), .DIA3(Data[39]), .DIA4(Data[40]), 
        .DIA5(Data[41]), .DIA6(Data[42]), .DIA7(Data[43]), .DIA8(Data[44]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_36), 
        .DOB1(mdout1_3_37), .DOB2(mdout1_3_38), .DOB3(mdout1_3_39), .DOB4(mdout1_3_40), 
        .DOB5(mdout1_3_41), .DOB6(mdout1_3_42), .DOB7(mdout1_3_43), .DOB8(mdout1_3_44), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49 (.DIA0(Data[45]), 
        .DIA1(Data[46]), .DIA2(Data[47]), .DIA3(Data[48]), .DIA4(Data[49]), 
        .DIA5(Data[50]), .DIA6(Data[51]), .DIA7(Data[52]), .DIA8(Data[53]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_45), 
        .DOB1(mdout1_3_46), .DOB2(mdout1_3_47), .DOB3(mdout1_3_48), .DOB4(mdout1_3_49), 
        .DOB5(mdout1_3_50), .DOB6(mdout1_3_51), .DOB7(mdout1_3_52), .DOB8(mdout1_3_53), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48 (.DIA0(Data[54]), 
        .DIA1(Data[55]), .DIA2(Data[56]), .DIA3(Data[57]), .DIA4(Data[58]), 
        .DIA5(Data[59]), .DIA6(Data[60]), .DIA7(Data[61]), .DIA8(Data[62]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_54), 
        .DOB1(mdout1_3_55), .DOB2(mdout1_3_56), .DOB3(mdout1_3_57), .DOB4(mdout1_3_58), 
        .DOB5(mdout1_3_59), .DOB6(mdout1_3_60), .DOB7(mdout1_3_61), .DOB8(mdout1_3_62), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47 (.DIA0(Data[63]), 
        .DIA1(Data[64]), .DIA2(Data[65]), .DIA3(Data[66]), .DIA4(Data[67]), 
        .DIA5(Data[68]), .DIA6(Data[69]), .DIA7(Data[70]), .DIA8(Data[71]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_63), 
        .DOB1(mdout1_3_64), .DOB2(mdout1_3_65), .DOB3(mdout1_3_66), .DOB4(mdout1_3_67), 
        .DOB5(mdout1_3_68), .DOB6(mdout1_3_69), .DOB7(mdout1_3_70), .DOB8(mdout1_3_71), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46 (.DIA0(Data[72]), 
        .DIA1(Data[73]), .DIA2(Data[74]), .DIA3(Data[75]), .DIA4(Data[76]), 
        .DIA5(Data[77]), .DIA6(Data[78]), .DIA7(Data[79]), .DIA8(Data[80]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_72), 
        .DOB1(mdout1_3_73), .DOB2(mdout1_3_74), .DOB3(mdout1_3_75), .DOB4(mdout1_3_76), 
        .DOB5(mdout1_3_77), .DOB6(mdout1_3_78), .DOB7(mdout1_3_79), .DOB8(mdout1_3_80), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45 (.DIA0(Data[81]), 
        .DIA1(Data[82]), .DIA2(Data[83]), .DIA3(Data[84]), .DIA4(Data[85]), 
        .DIA5(Data[86]), .DIA6(Data[87]), .DIA7(Data[88]), .DIA8(Data[89]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_81), 
        .DOB1(mdout1_3_82), .DOB2(mdout1_3_83), .DOB3(mdout1_3_84), .DOB4(mdout1_3_85), 
        .DOB5(mdout1_3_86), .DOB6(mdout1_3_87), .DOB7(mdout1_3_88), .DOB8(mdout1_3_89), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44.CSDECODE_B = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44.CSDECODE_A = "0b011" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44 (.DIA0(Data[90]), 
        .DIA1(Data[91]), .DIA2(Data[92]), .DIA3(Data[93]), .DIA4(Data[94]), 
        .DIA5(Data[95]), .DIA6(Data[96]), .DIA7(Data[97]), .DIA8(Data[98]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_3_90), 
        .DOB1(mdout1_3_91), .DOB2(mdout1_3_92), .DOB3(mdout1_3_93), .DOB4(mdout1_3_94), 
        .DOB5(mdout1_3_95), .DOB6(mdout1_3_96), .DOB7(mdout1_3_97), .DOB8(mdout1_3_98), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43 (.DIA0(Data[0]), 
        .DIA1(Data[1]), .DIA2(Data[2]), .DIA3(Data[3]), .DIA4(Data[4]), 
        .DIA5(Data[5]), .DIA6(Data[6]), .DIA7(Data[7]), .DIA8(Data[8]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_0), 
        .DOB1(mdout1_4_1), .DOB2(mdout1_4_2), .DOB3(mdout1_4_3), .DOB4(mdout1_4_4), 
        .DOB5(mdout1_4_5), .DOB6(mdout1_4_6), .DOB7(mdout1_4_7), .DOB8(mdout1_4_8), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42 (.DIA0(Data[9]), 
        .DIA1(Data[10]), .DIA2(Data[11]), .DIA3(Data[12]), .DIA4(Data[13]), 
        .DIA5(Data[14]), .DIA6(Data[15]), .DIA7(Data[16]), .DIA8(Data[17]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_9), 
        .DOB1(mdout1_4_10), .DOB2(mdout1_4_11), .DOB3(mdout1_4_12), .DOB4(mdout1_4_13), 
        .DOB5(mdout1_4_14), .DOB6(mdout1_4_15), .DOB7(mdout1_4_16), .DOB8(mdout1_4_17), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41 (.DIA0(Data[18]), 
        .DIA1(Data[19]), .DIA2(Data[20]), .DIA3(Data[21]), .DIA4(Data[22]), 
        .DIA5(Data[23]), .DIA6(Data[24]), .DIA7(Data[25]), .DIA8(Data[26]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_18), 
        .DOB1(mdout1_4_19), .DOB2(mdout1_4_20), .DOB3(mdout1_4_21), .DOB4(mdout1_4_22), 
        .DOB5(mdout1_4_23), .DOB6(mdout1_4_24), .DOB7(mdout1_4_25), .DOB8(mdout1_4_26), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40 (.DIA0(Data[27]), 
        .DIA1(Data[28]), .DIA2(Data[29]), .DIA3(Data[30]), .DIA4(Data[31]), 
        .DIA5(Data[32]), .DIA6(Data[33]), .DIA7(Data[34]), .DIA8(Data[35]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_27), 
        .DOB1(mdout1_4_28), .DOB2(mdout1_4_29), .DOB3(mdout1_4_30), .DOB4(mdout1_4_31), 
        .DOB5(mdout1_4_32), .DOB6(mdout1_4_33), .DOB7(mdout1_4_34), .DOB8(mdout1_4_35), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39 (.DIA0(Data[36]), 
        .DIA1(Data[37]), .DIA2(Data[38]), .DIA3(Data[39]), .DIA4(Data[40]), 
        .DIA5(Data[41]), .DIA6(Data[42]), .DIA7(Data[43]), .DIA8(Data[44]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_36), 
        .DOB1(mdout1_4_37), .DOB2(mdout1_4_38), .DOB3(mdout1_4_39), .DOB4(mdout1_4_40), 
        .DOB5(mdout1_4_41), .DOB6(mdout1_4_42), .DOB7(mdout1_4_43), .DOB8(mdout1_4_44), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38 (.DIA0(Data[45]), 
        .DIA1(Data[46]), .DIA2(Data[47]), .DIA3(Data[48]), .DIA4(Data[49]), 
        .DIA5(Data[50]), .DIA6(Data[51]), .DIA7(Data[52]), .DIA8(Data[53]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_45), 
        .DOB1(mdout1_4_46), .DOB2(mdout1_4_47), .DOB3(mdout1_4_48), .DOB4(mdout1_4_49), 
        .DOB5(mdout1_4_50), .DOB6(mdout1_4_51), .DOB7(mdout1_4_52), .DOB8(mdout1_4_53), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37 (.DIA0(Data[54]), 
        .DIA1(Data[55]), .DIA2(Data[56]), .DIA3(Data[57]), .DIA4(Data[58]), 
        .DIA5(Data[59]), .DIA6(Data[60]), .DIA7(Data[61]), .DIA8(Data[62]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_54), 
        .DOB1(mdout1_4_55), .DOB2(mdout1_4_56), .DOB3(mdout1_4_57), .DOB4(mdout1_4_58), 
        .DOB5(mdout1_4_59), .DOB6(mdout1_4_60), .DOB7(mdout1_4_61), .DOB8(mdout1_4_62), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36 (.DIA0(Data[63]), 
        .DIA1(Data[64]), .DIA2(Data[65]), .DIA3(Data[66]), .DIA4(Data[67]), 
        .DIA5(Data[68]), .DIA6(Data[69]), .DIA7(Data[70]), .DIA8(Data[71]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_63), 
        .DOB1(mdout1_4_64), .DOB2(mdout1_4_65), .DOB3(mdout1_4_66), .DOB4(mdout1_4_67), 
        .DOB5(mdout1_4_68), .DOB6(mdout1_4_69), .DOB7(mdout1_4_70), .DOB8(mdout1_4_71), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35 (.DIA0(Data[72]), 
        .DIA1(Data[73]), .DIA2(Data[74]), .DIA3(Data[75]), .DIA4(Data[76]), 
        .DIA5(Data[77]), .DIA6(Data[78]), .DIA7(Data[79]), .DIA8(Data[80]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_72), 
        .DOB1(mdout1_4_73), .DOB2(mdout1_4_74), .DOB3(mdout1_4_75), .DOB4(mdout1_4_76), 
        .DOB5(mdout1_4_77), .DOB6(mdout1_4_78), .DOB7(mdout1_4_79), .DOB8(mdout1_4_80), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34 (.DIA0(Data[81]), 
        .DIA1(Data[82]), .DIA2(Data[83]), .DIA3(Data[84]), .DIA4(Data[85]), 
        .DIA5(Data[86]), .DIA6(Data[87]), .DIA7(Data[88]), .DIA8(Data[89]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_81), 
        .DOB1(mdout1_4_82), .DOB2(mdout1_4_83), .DOB3(mdout1_4_84), .DOB4(mdout1_4_85), 
        .DOB5(mdout1_4_86), .DOB6(mdout1_4_87), .DOB7(mdout1_4_88), .DOB8(mdout1_4_89), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33.CSDECODE_B = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33.CSDECODE_A = "0b100" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33 (.DIA0(Data[90]), 
        .DIA1(Data[91]), .DIA2(Data[92]), .DIA3(Data[93]), .DIA4(Data[94]), 
        .DIA5(Data[95]), .DIA6(Data[96]), .DIA7(Data[97]), .DIA8(Data[98]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_4_90), 
        .DOB1(mdout1_4_91), .DOB2(mdout1_4_92), .DOB3(mdout1_4_93), .DOB4(mdout1_4_94), 
        .DOB5(mdout1_4_95), .DOB6(mdout1_4_96), .DOB7(mdout1_4_97), .DOB8(mdout1_4_98), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32 (.DIA0(Data[0]), 
        .DIA1(Data[1]), .DIA2(Data[2]), .DIA3(Data[3]), .DIA4(Data[4]), 
        .DIA5(Data[5]), .DIA6(Data[6]), .DIA7(Data[7]), .DIA8(Data[8]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_0), 
        .DOB1(mdout1_5_1), .DOB2(mdout1_5_2), .DOB3(mdout1_5_3), .DOB4(mdout1_5_4), 
        .DOB5(mdout1_5_5), .DOB6(mdout1_5_6), .DOB7(mdout1_5_7), .DOB8(mdout1_5_8), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31 (.DIA0(Data[9]), 
        .DIA1(Data[10]), .DIA2(Data[11]), .DIA3(Data[12]), .DIA4(Data[13]), 
        .DIA5(Data[14]), .DIA6(Data[15]), .DIA7(Data[16]), .DIA8(Data[17]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_9), 
        .DOB1(mdout1_5_10), .DOB2(mdout1_5_11), .DOB3(mdout1_5_12), .DOB4(mdout1_5_13), 
        .DOB5(mdout1_5_14), .DOB6(mdout1_5_15), .DOB7(mdout1_5_16), .DOB8(mdout1_5_17), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30 (.DIA0(Data[18]), 
        .DIA1(Data[19]), .DIA2(Data[20]), .DIA3(Data[21]), .DIA4(Data[22]), 
        .DIA5(Data[23]), .DIA6(Data[24]), .DIA7(Data[25]), .DIA8(Data[26]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_18), 
        .DOB1(mdout1_5_19), .DOB2(mdout1_5_20), .DOB3(mdout1_5_21), .DOB4(mdout1_5_22), 
        .DOB5(mdout1_5_23), .DOB6(mdout1_5_24), .DOB7(mdout1_5_25), .DOB8(mdout1_5_26), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29 (.DIA0(Data[27]), 
        .DIA1(Data[28]), .DIA2(Data[29]), .DIA3(Data[30]), .DIA4(Data[31]), 
        .DIA5(Data[32]), .DIA6(Data[33]), .DIA7(Data[34]), .DIA8(Data[35]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_27), 
        .DOB1(mdout1_5_28), .DOB2(mdout1_5_29), .DOB3(mdout1_5_30), .DOB4(mdout1_5_31), 
        .DOB5(mdout1_5_32), .DOB6(mdout1_5_33), .DOB7(mdout1_5_34), .DOB8(mdout1_5_35), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28 (.DIA0(Data[36]), 
        .DIA1(Data[37]), .DIA2(Data[38]), .DIA3(Data[39]), .DIA4(Data[40]), 
        .DIA5(Data[41]), .DIA6(Data[42]), .DIA7(Data[43]), .DIA8(Data[44]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_36), 
        .DOB1(mdout1_5_37), .DOB2(mdout1_5_38), .DOB3(mdout1_5_39), .DOB4(mdout1_5_40), 
        .DOB5(mdout1_5_41), .DOB6(mdout1_5_42), .DOB7(mdout1_5_43), .DOB8(mdout1_5_44), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27 (.DIA0(Data[45]), 
        .DIA1(Data[46]), .DIA2(Data[47]), .DIA3(Data[48]), .DIA4(Data[49]), 
        .DIA5(Data[50]), .DIA6(Data[51]), .DIA7(Data[52]), .DIA8(Data[53]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_45), 
        .DOB1(mdout1_5_46), .DOB2(mdout1_5_47), .DOB3(mdout1_5_48), .DOB4(mdout1_5_49), 
        .DOB5(mdout1_5_50), .DOB6(mdout1_5_51), .DOB7(mdout1_5_52), .DOB8(mdout1_5_53), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26 (.DIA0(Data[54]), 
        .DIA1(Data[55]), .DIA2(Data[56]), .DIA3(Data[57]), .DIA4(Data[58]), 
        .DIA5(Data[59]), .DIA6(Data[60]), .DIA7(Data[61]), .DIA8(Data[62]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_54), 
        .DOB1(mdout1_5_55), .DOB2(mdout1_5_56), .DOB3(mdout1_5_57), .DOB4(mdout1_5_58), 
        .DOB5(mdout1_5_59), .DOB6(mdout1_5_60), .DOB7(mdout1_5_61), .DOB8(mdout1_5_62), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25 (.DIA0(Data[63]), 
        .DIA1(Data[64]), .DIA2(Data[65]), .DIA3(Data[66]), .DIA4(Data[67]), 
        .DIA5(Data[68]), .DIA6(Data[69]), .DIA7(Data[70]), .DIA8(Data[71]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_63), 
        .DOB1(mdout1_5_64), .DOB2(mdout1_5_65), .DOB3(mdout1_5_66), .DOB4(mdout1_5_67), 
        .DOB5(mdout1_5_68), .DOB6(mdout1_5_69), .DOB7(mdout1_5_70), .DOB8(mdout1_5_71), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24 (.DIA0(Data[72]), 
        .DIA1(Data[73]), .DIA2(Data[74]), .DIA3(Data[75]), .DIA4(Data[76]), 
        .DIA5(Data[77]), .DIA6(Data[78]), .DIA7(Data[79]), .DIA8(Data[80]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_72), 
        .DOB1(mdout1_5_73), .DOB2(mdout1_5_74), .DOB3(mdout1_5_75), .DOB4(mdout1_5_76), 
        .DOB5(mdout1_5_77), .DOB6(mdout1_5_78), .DOB7(mdout1_5_79), .DOB8(mdout1_5_80), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23 (.DIA0(Data[81]), 
        .DIA1(Data[82]), .DIA2(Data[83]), .DIA3(Data[84]), .DIA4(Data[85]), 
        .DIA5(Data[86]), .DIA6(Data[87]), .DIA7(Data[88]), .DIA8(Data[89]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_81), 
        .DOB1(mdout1_5_82), .DOB2(mdout1_5_83), .DOB3(mdout1_5_84), .DOB4(mdout1_5_85), 
        .DOB5(mdout1_5_86), .DOB6(mdout1_5_87), .DOB7(mdout1_5_88), .DOB8(mdout1_5_89), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22.CSDECODE_B = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22.CSDECODE_A = "0b101" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22 (.DIA0(Data[90]), 
        .DIA1(Data[91]), .DIA2(Data[92]), .DIA3(Data[93]), .DIA4(Data[94]), 
        .DIA5(Data[95]), .DIA6(Data[96]), .DIA7(Data[97]), .DIA8(Data[98]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_5_90), 
        .DOB1(mdout1_5_91), .DOB2(mdout1_5_92), .DOB3(mdout1_5_93), .DOB4(mdout1_5_94), 
        .DOB5(mdout1_5_95), .DOB6(mdout1_5_96), .DOB7(mdout1_5_97), .DOB8(mdout1_5_98), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21 (.DIA0(Data[0]), 
        .DIA1(Data[1]), .DIA2(Data[2]), .DIA3(Data[3]), .DIA4(Data[4]), 
        .DIA5(Data[5]), .DIA6(Data[6]), .DIA7(Data[7]), .DIA8(Data[8]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_0), 
        .DOB1(mdout1_6_1), .DOB2(mdout1_6_2), .DOB3(mdout1_6_3), .DOB4(mdout1_6_4), 
        .DOB5(mdout1_6_5), .DOB6(mdout1_6_6), .DOB7(mdout1_6_7), .DOB8(mdout1_6_8), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20 (.DIA0(Data[9]), 
        .DIA1(Data[10]), .DIA2(Data[11]), .DIA3(Data[12]), .DIA4(Data[13]), 
        .DIA5(Data[14]), .DIA6(Data[15]), .DIA7(Data[16]), .DIA8(Data[17]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_9), 
        .DOB1(mdout1_6_10), .DOB2(mdout1_6_11), .DOB3(mdout1_6_12), .DOB4(mdout1_6_13), 
        .DOB5(mdout1_6_14), .DOB6(mdout1_6_15), .DOB7(mdout1_6_16), .DOB8(mdout1_6_17), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19 (.DIA0(Data[18]), 
        .DIA1(Data[19]), .DIA2(Data[20]), .DIA3(Data[21]), .DIA4(Data[22]), 
        .DIA5(Data[23]), .DIA6(Data[24]), .DIA7(Data[25]), .DIA8(Data[26]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_18), 
        .DOB1(mdout1_6_19), .DOB2(mdout1_6_20), .DOB3(mdout1_6_21), .DOB4(mdout1_6_22), 
        .DOB5(mdout1_6_23), .DOB6(mdout1_6_24), .DOB7(mdout1_6_25), .DOB8(mdout1_6_26), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18 (.DIA0(Data[27]), 
        .DIA1(Data[28]), .DIA2(Data[29]), .DIA3(Data[30]), .DIA4(Data[31]), 
        .DIA5(Data[32]), .DIA6(Data[33]), .DIA7(Data[34]), .DIA8(Data[35]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_27), 
        .DOB1(mdout1_6_28), .DOB2(mdout1_6_29), .DOB3(mdout1_6_30), .DOB4(mdout1_6_31), 
        .DOB5(mdout1_6_32), .DOB6(mdout1_6_33), .DOB7(mdout1_6_34), .DOB8(mdout1_6_35), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17 (.DIA0(Data[36]), 
        .DIA1(Data[37]), .DIA2(Data[38]), .DIA3(Data[39]), .DIA4(Data[40]), 
        .DIA5(Data[41]), .DIA6(Data[42]), .DIA7(Data[43]), .DIA8(Data[44]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_36), 
        .DOB1(mdout1_6_37), .DOB2(mdout1_6_38), .DOB3(mdout1_6_39), .DOB4(mdout1_6_40), 
        .DOB5(mdout1_6_41), .DOB6(mdout1_6_42), .DOB7(mdout1_6_43), .DOB8(mdout1_6_44), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16 (.DIA0(Data[45]), 
        .DIA1(Data[46]), .DIA2(Data[47]), .DIA3(Data[48]), .DIA4(Data[49]), 
        .DIA5(Data[50]), .DIA6(Data[51]), .DIA7(Data[52]), .DIA8(Data[53]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_45), 
        .DOB1(mdout1_6_46), .DOB2(mdout1_6_47), .DOB3(mdout1_6_48), .DOB4(mdout1_6_49), 
        .DOB5(mdout1_6_50), .DOB6(mdout1_6_51), .DOB7(mdout1_6_52), .DOB8(mdout1_6_53), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15 (.DIA0(Data[54]), 
        .DIA1(Data[55]), .DIA2(Data[56]), .DIA3(Data[57]), .DIA4(Data[58]), 
        .DIA5(Data[59]), .DIA6(Data[60]), .DIA7(Data[61]), .DIA8(Data[62]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_54), 
        .DOB1(mdout1_6_55), .DOB2(mdout1_6_56), .DOB3(mdout1_6_57), .DOB4(mdout1_6_58), 
        .DOB5(mdout1_6_59), .DOB6(mdout1_6_60), .DOB7(mdout1_6_61), .DOB8(mdout1_6_62), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14 (.DIA0(Data[63]), 
        .DIA1(Data[64]), .DIA2(Data[65]), .DIA3(Data[66]), .DIA4(Data[67]), 
        .DIA5(Data[68]), .DIA6(Data[69]), .DIA7(Data[70]), .DIA8(Data[71]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_63), 
        .DOB1(mdout1_6_64), .DOB2(mdout1_6_65), .DOB3(mdout1_6_66), .DOB4(mdout1_6_67), 
        .DOB5(mdout1_6_68), .DOB6(mdout1_6_69), .DOB7(mdout1_6_70), .DOB8(mdout1_6_71), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13 (.DIA0(Data[72]), 
        .DIA1(Data[73]), .DIA2(Data[74]), .DIA3(Data[75]), .DIA4(Data[76]), 
        .DIA5(Data[77]), .DIA6(Data[78]), .DIA7(Data[79]), .DIA8(Data[80]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_72), 
        .DOB1(mdout1_6_73), .DOB2(mdout1_6_74), .DOB3(mdout1_6_75), .DOB4(mdout1_6_76), 
        .DOB5(mdout1_6_77), .DOB6(mdout1_6_78), .DOB7(mdout1_6_79), .DOB8(mdout1_6_80), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12 (.DIA0(Data[81]), 
        .DIA1(Data[82]), .DIA2(Data[83]), .DIA3(Data[84]), .DIA4(Data[85]), 
        .DIA5(Data[86]), .DIA6(Data[87]), .DIA7(Data[88]), .DIA8(Data[89]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_81), 
        .DOB1(mdout1_6_82), .DOB2(mdout1_6_83), .DOB3(mdout1_6_84), .DOB4(mdout1_6_85), 
        .DOB5(mdout1_6_86), .DOB6(mdout1_6_87), .DOB7(mdout1_6_88), .DOB8(mdout1_6_89), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11.CSDECODE_B = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11.CSDECODE_A = "0b110" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11 (.DIA0(Data[90]), 
        .DIA1(Data[91]), .DIA2(Data[92]), .DIA3(Data[93]), .DIA4(Data[94]), 
        .DIA5(Data[95]), .DIA6(Data[96]), .DIA7(Data[97]), .DIA8(Data[98]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_6_90), 
        .DOB1(mdout1_6_91), .DOB2(mdout1_6_92), .DOB3(mdout1_6_93), .DOB4(mdout1_6_94), 
        .DOB5(mdout1_6_95), .DOB6(mdout1_6_96), .DOB7(mdout1_6_97), .DOB8(mdout1_6_98), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10 (.DIA0(Data[0]), 
        .DIA1(Data[1]), .DIA2(Data[2]), .DIA3(Data[3]), .DIA4(Data[4]), 
        .DIA5(Data[5]), .DIA6(Data[6]), .DIA7(Data[7]), .DIA8(Data[8]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_0), 
        .DOB1(mdout1_7_1), .DOB2(mdout1_7_2), .DOB3(mdout1_7_3), .DOB4(mdout1_7_4), 
        .DOB5(mdout1_7_5), .DOB6(mdout1_7_6), .DOB7(mdout1_7_7), .DOB8(mdout1_7_8), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9 (.DIA0(Data[9]), 
        .DIA1(Data[10]), .DIA2(Data[11]), .DIA3(Data[12]), .DIA4(Data[13]), 
        .DIA5(Data[14]), .DIA6(Data[15]), .DIA7(Data[16]), .DIA8(Data[17]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_9), 
        .DOB1(mdout1_7_10), .DOB2(mdout1_7_11), .DOB3(mdout1_7_12), .DOB4(mdout1_7_13), 
        .DOB5(mdout1_7_14), .DOB6(mdout1_7_15), .DOB7(mdout1_7_16), .DOB8(mdout1_7_17), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8 (.DIA0(Data[18]), 
        .DIA1(Data[19]), .DIA2(Data[20]), .DIA3(Data[21]), .DIA4(Data[22]), 
        .DIA5(Data[23]), .DIA6(Data[24]), .DIA7(Data[25]), .DIA8(Data[26]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_18), 
        .DOB1(mdout1_7_19), .DOB2(mdout1_7_20), .DOB3(mdout1_7_21), .DOB4(mdout1_7_22), 
        .DOB5(mdout1_7_23), .DOB6(mdout1_7_24), .DOB7(mdout1_7_25), .DOB8(mdout1_7_26), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7 (.DIA0(Data[27]), 
        .DIA1(Data[28]), .DIA2(Data[29]), .DIA3(Data[30]), .DIA4(Data[31]), 
        .DIA5(Data[32]), .DIA6(Data[33]), .DIA7(Data[34]), .DIA8(Data[35]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_27), 
        .DOB1(mdout1_7_28), .DOB2(mdout1_7_29), .DOB3(mdout1_7_30), .DOB4(mdout1_7_31), 
        .DOB5(mdout1_7_32), .DOB6(mdout1_7_33), .DOB7(mdout1_7_34), .DOB8(mdout1_7_35), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6 (.DIA0(Data[36]), 
        .DIA1(Data[37]), .DIA2(Data[38]), .DIA3(Data[39]), .DIA4(Data[40]), 
        .DIA5(Data[41]), .DIA6(Data[42]), .DIA7(Data[43]), .DIA8(Data[44]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_36), 
        .DOB1(mdout1_7_37), .DOB2(mdout1_7_38), .DOB3(mdout1_7_39), .DOB4(mdout1_7_40), 
        .DOB5(mdout1_7_41), .DOB6(mdout1_7_42), .DOB7(mdout1_7_43), .DOB8(mdout1_7_44), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5 (.DIA0(Data[45]), 
        .DIA1(Data[46]), .DIA2(Data[47]), .DIA3(Data[48]), .DIA4(Data[49]), 
        .DIA5(Data[50]), .DIA6(Data[51]), .DIA7(Data[52]), .DIA8(Data[53]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_45), 
        .DOB1(mdout1_7_46), .DOB2(mdout1_7_47), .DOB3(mdout1_7_48), .DOB4(mdout1_7_49), 
        .DOB5(mdout1_7_50), .DOB6(mdout1_7_51), .DOB7(mdout1_7_52), .DOB8(mdout1_7_53), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4 (.DIA0(Data[54]), 
        .DIA1(Data[55]), .DIA2(Data[56]), .DIA3(Data[57]), .DIA4(Data[58]), 
        .DIA5(Data[59]), .DIA6(Data[60]), .DIA7(Data[61]), .DIA8(Data[62]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_54), 
        .DOB1(mdout1_7_55), .DOB2(mdout1_7_56), .DOB3(mdout1_7_57), .DOB4(mdout1_7_58), 
        .DOB5(mdout1_7_59), .DOB6(mdout1_7_60), .DOB7(mdout1_7_61), .DOB8(mdout1_7_62), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3 (.DIA0(Data[63]), 
        .DIA1(Data[64]), .DIA2(Data[65]), .DIA3(Data[66]), .DIA4(Data[67]), 
        .DIA5(Data[68]), .DIA6(Data[69]), .DIA7(Data[70]), .DIA8(Data[71]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_63), 
        .DOB1(mdout1_7_64), .DOB2(mdout1_7_65), .DOB3(mdout1_7_66), .DOB4(mdout1_7_67), 
        .DOB5(mdout1_7_68), .DOB6(mdout1_7_69), .DOB7(mdout1_7_70), .DOB8(mdout1_7_71), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2 (.DIA0(Data[72]), 
        .DIA1(Data[73]), .DIA2(Data[74]), .DIA3(Data[75]), .DIA4(Data[76]), 
        .DIA5(Data[77]), .DIA6(Data[78]), .DIA7(Data[79]), .DIA8(Data[80]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_72), 
        .DOB1(mdout1_7_73), .DOB2(mdout1_7_74), .DOB3(mdout1_7_75), .DOB4(mdout1_7_76), 
        .DOB5(mdout1_7_77), .DOB6(mdout1_7_78), .DOB7(mdout1_7_79), .DOB8(mdout1_7_80), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1 (.DIA0(Data[81]), 
        .DIA1(Data[82]), .DIA2(Data[83]), .DIA3(Data[84]), .DIA4(Data[85]), 
        .DIA5(Data[86]), .DIA6(Data[87]), .DIA7(Data[88]), .DIA8(Data[89]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_81), 
        .DOB1(mdout1_7_82), .DOB2(mdout1_7_83), .DOB3(mdout1_7_84), .DOB4(mdout1_7_85), 
        .DOB5(mdout1_7_86), .DOB6(mdout1_7_87), .DOB7(mdout1_7_88), .DOB8(mdout1_7_89), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0.CSDECODE_B = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0.CSDECODE_A = "0b111" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0.GSR = "DISABLED" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0.DATA_WIDTH_A = 9 ;
    DP16KC pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0 (.DIA0(Data[90]), 
        .DIA1(Data[91]), .DIA2(Data[92]), .DIA3(Data[93]), .DIA4(Data[94]), 
        .DIA5(Data[95]), .DIA6(Data[96]), .DIA7(Data[97]), .DIA8(Data[98]), 
        .DIA9(scuba_vlo), .DIA10(scuba_vlo), .DIA11(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA13(scuba_vlo), .DIA14(scuba_vlo), .DIA15(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA17(scuba_vlo), .ADA0(scuba_vlo), .ADA1(scuba_vlo), .ADA2(scuba_vlo), 
        .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), 
        .ADA7(WrAddress[4]), .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
        .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
        .CEA(WrClockEn), .CLKA(WrClock), .OCEA(WrClockEn), .WEA(WE), .CSA0(WrAddress[11]), 
        .CSA1(WrAddress[12]), .CSA2(WrAddress[13]), .RSTA(Reset), .DIB0(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), 
        .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), 
        .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
        .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
        .CEB(RdClockEn), .CLKB(RdClock), .OCEB(RdClockEn), .WEB(scuba_vlo), 
        .CSB0(RdAddress[11]), .CSB1(RdAddress[12]), .CSB2(RdAddress[13]), 
        .RSTB(Reset), .DOA0(), .DOA1(), .DOA2(), .DOA3(), .DOA4(), .DOA5(), 
        .DOA6(), .DOA7(), .DOA8(), .DOA9(), .DOA10(), .DOA11(), .DOA12(), 
        .DOA13(), .DOA14(), .DOA15(), .DOA16(), .DOA17(), .DOB0(mdout1_7_90), 
        .DOB1(mdout1_7_91), .DOB2(mdout1_7_92), .DOB3(mdout1_7_93), .DOB4(mdout1_7_94), 
        .DOB5(mdout1_7_95), .DOB6(mdout1_7_96), .DOB7(mdout1_7_97), .DOB8(mdout1_7_98), 
        .DOB9(), .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), 
        .DOB16(), .DOB17())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B" */
             /* synthesis MEM_INIT_FILE="" */
             /* synthesis RESETMODE="SYNC" */;

    FD1P3DX FF_5 (.D(RdAddress[11]), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr11_ff))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_4 (.D(RdAddress[12]), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr12_ff))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_3 (.D(RdAddress[13]), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr13_ff))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_2 (.D(raddr11_ff), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr11_ff2))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_1 (.D(raddr12_ff), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr12_ff2))
             /* synthesis GSR="ENABLED" */;

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    FD1P3DX FF_0 (.D(raddr13_ff), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr13_ff2))
             /* synthesis GSR="ENABLED" */;

    MUX81 mux_98 (.D0(mdout1_0_0), .D1(mdout1_1_0), .D2(mdout1_2_0), .D3(mdout1_3_0), 
        .D4(mdout1_4_0), .D5(mdout1_5_0), .D6(mdout1_6_0), .D7(mdout1_7_0), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[0]));

    MUX81 mux_97 (.D0(mdout1_0_1), .D1(mdout1_1_1), .D2(mdout1_2_1), .D3(mdout1_3_1), 
        .D4(mdout1_4_1), .D5(mdout1_5_1), .D6(mdout1_6_1), .D7(mdout1_7_1), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[1]));

    MUX81 mux_96 (.D0(mdout1_0_2), .D1(mdout1_1_2), .D2(mdout1_2_2), .D3(mdout1_3_2), 
        .D4(mdout1_4_2), .D5(mdout1_5_2), .D6(mdout1_6_2), .D7(mdout1_7_2), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[2]));

    MUX81 mux_95 (.D0(mdout1_0_3), .D1(mdout1_1_3), .D2(mdout1_2_3), .D3(mdout1_3_3), 
        .D4(mdout1_4_3), .D5(mdout1_5_3), .D6(mdout1_6_3), .D7(mdout1_7_3), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[3]));

    MUX81 mux_94 (.D0(mdout1_0_4), .D1(mdout1_1_4), .D2(mdout1_2_4), .D3(mdout1_3_4), 
        .D4(mdout1_4_4), .D5(mdout1_5_4), .D6(mdout1_6_4), .D7(mdout1_7_4), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[4]));

    MUX81 mux_93 (.D0(mdout1_0_5), .D1(mdout1_1_5), .D2(mdout1_2_5), .D3(mdout1_3_5), 
        .D4(mdout1_4_5), .D5(mdout1_5_5), .D6(mdout1_6_5), .D7(mdout1_7_5), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[5]));

    MUX81 mux_92 (.D0(mdout1_0_6), .D1(mdout1_1_6), .D2(mdout1_2_6), .D3(mdout1_3_6), 
        .D4(mdout1_4_6), .D5(mdout1_5_6), .D6(mdout1_6_6), .D7(mdout1_7_6), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[6]));

    MUX81 mux_91 (.D0(mdout1_0_7), .D1(mdout1_1_7), .D2(mdout1_2_7), .D3(mdout1_3_7), 
        .D4(mdout1_4_7), .D5(mdout1_5_7), .D6(mdout1_6_7), .D7(mdout1_7_7), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[7]));

    MUX81 mux_90 (.D0(mdout1_0_8), .D1(mdout1_1_8), .D2(mdout1_2_8), .D3(mdout1_3_8), 
        .D4(mdout1_4_8), .D5(mdout1_5_8), .D6(mdout1_6_8), .D7(mdout1_7_8), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[8]));

    MUX81 mux_89 (.D0(mdout1_0_9), .D1(mdout1_1_9), .D2(mdout1_2_9), .D3(mdout1_3_9), 
        .D4(mdout1_4_9), .D5(mdout1_5_9), .D6(mdout1_6_9), .D7(mdout1_7_9), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[9]));

    MUX81 mux_88 (.D0(mdout1_0_10), .D1(mdout1_1_10), .D2(mdout1_2_10), 
        .D3(mdout1_3_10), .D4(mdout1_4_10), .D5(mdout1_5_10), .D6(mdout1_6_10), 
        .D7(mdout1_7_10), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[10]));

    MUX81 mux_87 (.D0(mdout1_0_11), .D1(mdout1_1_11), .D2(mdout1_2_11), 
        .D3(mdout1_3_11), .D4(mdout1_4_11), .D5(mdout1_5_11), .D6(mdout1_6_11), 
        .D7(mdout1_7_11), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[11]));

    MUX81 mux_86 (.D0(mdout1_0_12), .D1(mdout1_1_12), .D2(mdout1_2_12), 
        .D3(mdout1_3_12), .D4(mdout1_4_12), .D5(mdout1_5_12), .D6(mdout1_6_12), 
        .D7(mdout1_7_12), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[12]));

    MUX81 mux_85 (.D0(mdout1_0_13), .D1(mdout1_1_13), .D2(mdout1_2_13), 
        .D3(mdout1_3_13), .D4(mdout1_4_13), .D5(mdout1_5_13), .D6(mdout1_6_13), 
        .D7(mdout1_7_13), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[13]));

    MUX81 mux_84 (.D0(mdout1_0_14), .D1(mdout1_1_14), .D2(mdout1_2_14), 
        .D3(mdout1_3_14), .D4(mdout1_4_14), .D5(mdout1_5_14), .D6(mdout1_6_14), 
        .D7(mdout1_7_14), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[14]));

    MUX81 mux_83 (.D0(mdout1_0_15), .D1(mdout1_1_15), .D2(mdout1_2_15), 
        .D3(mdout1_3_15), .D4(mdout1_4_15), .D5(mdout1_5_15), .D6(mdout1_6_15), 
        .D7(mdout1_7_15), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[15]));

    MUX81 mux_82 (.D0(mdout1_0_16), .D1(mdout1_1_16), .D2(mdout1_2_16), 
        .D3(mdout1_3_16), .D4(mdout1_4_16), .D5(mdout1_5_16), .D6(mdout1_6_16), 
        .D7(mdout1_7_16), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[16]));

    MUX81 mux_81 (.D0(mdout1_0_17), .D1(mdout1_1_17), .D2(mdout1_2_17), 
        .D3(mdout1_3_17), .D4(mdout1_4_17), .D5(mdout1_5_17), .D6(mdout1_6_17), 
        .D7(mdout1_7_17), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[17]));

    MUX81 mux_80 (.D0(mdout1_0_18), .D1(mdout1_1_18), .D2(mdout1_2_18), 
        .D3(mdout1_3_18), .D4(mdout1_4_18), .D5(mdout1_5_18), .D6(mdout1_6_18), 
        .D7(mdout1_7_18), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[18]));

    MUX81 mux_79 (.D0(mdout1_0_19), .D1(mdout1_1_19), .D2(mdout1_2_19), 
        .D3(mdout1_3_19), .D4(mdout1_4_19), .D5(mdout1_5_19), .D6(mdout1_6_19), 
        .D7(mdout1_7_19), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[19]));

    MUX81 mux_78 (.D0(mdout1_0_20), .D1(mdout1_1_20), .D2(mdout1_2_20), 
        .D3(mdout1_3_20), .D4(mdout1_4_20), .D5(mdout1_5_20), .D6(mdout1_6_20), 
        .D7(mdout1_7_20), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[20]));

    MUX81 mux_77 (.D0(mdout1_0_21), .D1(mdout1_1_21), .D2(mdout1_2_21), 
        .D3(mdout1_3_21), .D4(mdout1_4_21), .D5(mdout1_5_21), .D6(mdout1_6_21), 
        .D7(mdout1_7_21), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[21]));

    MUX81 mux_76 (.D0(mdout1_0_22), .D1(mdout1_1_22), .D2(mdout1_2_22), 
        .D3(mdout1_3_22), .D4(mdout1_4_22), .D5(mdout1_5_22), .D6(mdout1_6_22), 
        .D7(mdout1_7_22), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[22]));

    MUX81 mux_75 (.D0(mdout1_0_23), .D1(mdout1_1_23), .D2(mdout1_2_23), 
        .D3(mdout1_3_23), .D4(mdout1_4_23), .D5(mdout1_5_23), .D6(mdout1_6_23), 
        .D7(mdout1_7_23), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[23]));

    MUX81 mux_74 (.D0(mdout1_0_24), .D1(mdout1_1_24), .D2(mdout1_2_24), 
        .D3(mdout1_3_24), .D4(mdout1_4_24), .D5(mdout1_5_24), .D6(mdout1_6_24), 
        .D7(mdout1_7_24), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[24]));

    MUX81 mux_73 (.D0(mdout1_0_25), .D1(mdout1_1_25), .D2(mdout1_2_25), 
        .D3(mdout1_3_25), .D4(mdout1_4_25), .D5(mdout1_5_25), .D6(mdout1_6_25), 
        .D7(mdout1_7_25), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[25]));

    MUX81 mux_72 (.D0(mdout1_0_26), .D1(mdout1_1_26), .D2(mdout1_2_26), 
        .D3(mdout1_3_26), .D4(mdout1_4_26), .D5(mdout1_5_26), .D6(mdout1_6_26), 
        .D7(mdout1_7_26), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[26]));

    MUX81 mux_71 (.D0(mdout1_0_27), .D1(mdout1_1_27), .D2(mdout1_2_27), 
        .D3(mdout1_3_27), .D4(mdout1_4_27), .D5(mdout1_5_27), .D6(mdout1_6_27), 
        .D7(mdout1_7_27), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[27]));

    MUX81 mux_70 (.D0(mdout1_0_28), .D1(mdout1_1_28), .D2(mdout1_2_28), 
        .D3(mdout1_3_28), .D4(mdout1_4_28), .D5(mdout1_5_28), .D6(mdout1_6_28), 
        .D7(mdout1_7_28), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[28]));

    MUX81 mux_69 (.D0(mdout1_0_29), .D1(mdout1_1_29), .D2(mdout1_2_29), 
        .D3(mdout1_3_29), .D4(mdout1_4_29), .D5(mdout1_5_29), .D6(mdout1_6_29), 
        .D7(mdout1_7_29), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[29]));

    MUX81 mux_68 (.D0(mdout1_0_30), .D1(mdout1_1_30), .D2(mdout1_2_30), 
        .D3(mdout1_3_30), .D4(mdout1_4_30), .D5(mdout1_5_30), .D6(mdout1_6_30), 
        .D7(mdout1_7_30), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[30]));

    MUX81 mux_67 (.D0(mdout1_0_31), .D1(mdout1_1_31), .D2(mdout1_2_31), 
        .D3(mdout1_3_31), .D4(mdout1_4_31), .D5(mdout1_5_31), .D6(mdout1_6_31), 
        .D7(mdout1_7_31), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[31]));

    MUX81 mux_66 (.D0(mdout1_0_32), .D1(mdout1_1_32), .D2(mdout1_2_32), 
        .D3(mdout1_3_32), .D4(mdout1_4_32), .D5(mdout1_5_32), .D6(mdout1_6_32), 
        .D7(mdout1_7_32), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[32]));

    MUX81 mux_65 (.D0(mdout1_0_33), .D1(mdout1_1_33), .D2(mdout1_2_33), 
        .D3(mdout1_3_33), .D4(mdout1_4_33), .D5(mdout1_5_33), .D6(mdout1_6_33), 
        .D7(mdout1_7_33), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[33]));

    MUX81 mux_64 (.D0(mdout1_0_34), .D1(mdout1_1_34), .D2(mdout1_2_34), 
        .D3(mdout1_3_34), .D4(mdout1_4_34), .D5(mdout1_5_34), .D6(mdout1_6_34), 
        .D7(mdout1_7_34), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[34]));

    MUX81 mux_63 (.D0(mdout1_0_35), .D1(mdout1_1_35), .D2(mdout1_2_35), 
        .D3(mdout1_3_35), .D4(mdout1_4_35), .D5(mdout1_5_35), .D6(mdout1_6_35), 
        .D7(mdout1_7_35), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[35]));

    MUX81 mux_62 (.D0(mdout1_0_36), .D1(mdout1_1_36), .D2(mdout1_2_36), 
        .D3(mdout1_3_36), .D4(mdout1_4_36), .D5(mdout1_5_36), .D6(mdout1_6_36), 
        .D7(mdout1_7_36), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[36]));

    MUX81 mux_61 (.D0(mdout1_0_37), .D1(mdout1_1_37), .D2(mdout1_2_37), 
        .D3(mdout1_3_37), .D4(mdout1_4_37), .D5(mdout1_5_37), .D6(mdout1_6_37), 
        .D7(mdout1_7_37), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[37]));

    MUX81 mux_60 (.D0(mdout1_0_38), .D1(mdout1_1_38), .D2(mdout1_2_38), 
        .D3(mdout1_3_38), .D4(mdout1_4_38), .D5(mdout1_5_38), .D6(mdout1_6_38), 
        .D7(mdout1_7_38), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[38]));

    MUX81 mux_59 (.D0(mdout1_0_39), .D1(mdout1_1_39), .D2(mdout1_2_39), 
        .D3(mdout1_3_39), .D4(mdout1_4_39), .D5(mdout1_5_39), .D6(mdout1_6_39), 
        .D7(mdout1_7_39), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[39]));

    MUX81 mux_58 (.D0(mdout1_0_40), .D1(mdout1_1_40), .D2(mdout1_2_40), 
        .D3(mdout1_3_40), .D4(mdout1_4_40), .D5(mdout1_5_40), .D6(mdout1_6_40), 
        .D7(mdout1_7_40), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[40]));

    MUX81 mux_57 (.D0(mdout1_0_41), .D1(mdout1_1_41), .D2(mdout1_2_41), 
        .D3(mdout1_3_41), .D4(mdout1_4_41), .D5(mdout1_5_41), .D6(mdout1_6_41), 
        .D7(mdout1_7_41), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[41]));

    MUX81 mux_56 (.D0(mdout1_0_42), .D1(mdout1_1_42), .D2(mdout1_2_42), 
        .D3(mdout1_3_42), .D4(mdout1_4_42), .D5(mdout1_5_42), .D6(mdout1_6_42), 
        .D7(mdout1_7_42), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[42]));

    MUX81 mux_55 (.D0(mdout1_0_43), .D1(mdout1_1_43), .D2(mdout1_2_43), 
        .D3(mdout1_3_43), .D4(mdout1_4_43), .D5(mdout1_5_43), .D6(mdout1_6_43), 
        .D7(mdout1_7_43), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[43]));

    MUX81 mux_54 (.D0(mdout1_0_44), .D1(mdout1_1_44), .D2(mdout1_2_44), 
        .D3(mdout1_3_44), .D4(mdout1_4_44), .D5(mdout1_5_44), .D6(mdout1_6_44), 
        .D7(mdout1_7_44), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[44]));

    MUX81 mux_53 (.D0(mdout1_0_45), .D1(mdout1_1_45), .D2(mdout1_2_45), 
        .D3(mdout1_3_45), .D4(mdout1_4_45), .D5(mdout1_5_45), .D6(mdout1_6_45), 
        .D7(mdout1_7_45), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[45]));

    MUX81 mux_52 (.D0(mdout1_0_46), .D1(mdout1_1_46), .D2(mdout1_2_46), 
        .D3(mdout1_3_46), .D4(mdout1_4_46), .D5(mdout1_5_46), .D6(mdout1_6_46), 
        .D7(mdout1_7_46), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[46]));

    MUX81 mux_51 (.D0(mdout1_0_47), .D1(mdout1_1_47), .D2(mdout1_2_47), 
        .D3(mdout1_3_47), .D4(mdout1_4_47), .D5(mdout1_5_47), .D6(mdout1_6_47), 
        .D7(mdout1_7_47), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[47]));

    MUX81 mux_50 (.D0(mdout1_0_48), .D1(mdout1_1_48), .D2(mdout1_2_48), 
        .D3(mdout1_3_48), .D4(mdout1_4_48), .D5(mdout1_5_48), .D6(mdout1_6_48), 
        .D7(mdout1_7_48), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[48]));

    MUX81 mux_49 (.D0(mdout1_0_49), .D1(mdout1_1_49), .D2(mdout1_2_49), 
        .D3(mdout1_3_49), .D4(mdout1_4_49), .D5(mdout1_5_49), .D6(mdout1_6_49), 
        .D7(mdout1_7_49), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[49]));

    MUX81 mux_48 (.D0(mdout1_0_50), .D1(mdout1_1_50), .D2(mdout1_2_50), 
        .D3(mdout1_3_50), .D4(mdout1_4_50), .D5(mdout1_5_50), .D6(mdout1_6_50), 
        .D7(mdout1_7_50), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[50]));

    MUX81 mux_47 (.D0(mdout1_0_51), .D1(mdout1_1_51), .D2(mdout1_2_51), 
        .D3(mdout1_3_51), .D4(mdout1_4_51), .D5(mdout1_5_51), .D6(mdout1_6_51), 
        .D7(mdout1_7_51), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[51]));

    MUX81 mux_46 (.D0(mdout1_0_52), .D1(mdout1_1_52), .D2(mdout1_2_52), 
        .D3(mdout1_3_52), .D4(mdout1_4_52), .D5(mdout1_5_52), .D6(mdout1_6_52), 
        .D7(mdout1_7_52), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[52]));

    MUX81 mux_45 (.D0(mdout1_0_53), .D1(mdout1_1_53), .D2(mdout1_2_53), 
        .D3(mdout1_3_53), .D4(mdout1_4_53), .D5(mdout1_5_53), .D6(mdout1_6_53), 
        .D7(mdout1_7_53), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[53]));

    MUX81 mux_44 (.D0(mdout1_0_54), .D1(mdout1_1_54), .D2(mdout1_2_54), 
        .D3(mdout1_3_54), .D4(mdout1_4_54), .D5(mdout1_5_54), .D6(mdout1_6_54), 
        .D7(mdout1_7_54), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[54]));

    MUX81 mux_43 (.D0(mdout1_0_55), .D1(mdout1_1_55), .D2(mdout1_2_55), 
        .D3(mdout1_3_55), .D4(mdout1_4_55), .D5(mdout1_5_55), .D6(mdout1_6_55), 
        .D7(mdout1_7_55), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[55]));

    MUX81 mux_42 (.D0(mdout1_0_56), .D1(mdout1_1_56), .D2(mdout1_2_56), 
        .D3(mdout1_3_56), .D4(mdout1_4_56), .D5(mdout1_5_56), .D6(mdout1_6_56), 
        .D7(mdout1_7_56), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[56]));

    MUX81 mux_41 (.D0(mdout1_0_57), .D1(mdout1_1_57), .D2(mdout1_2_57), 
        .D3(mdout1_3_57), .D4(mdout1_4_57), .D5(mdout1_5_57), .D6(mdout1_6_57), 
        .D7(mdout1_7_57), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[57]));

    MUX81 mux_40 (.D0(mdout1_0_58), .D1(mdout1_1_58), .D2(mdout1_2_58), 
        .D3(mdout1_3_58), .D4(mdout1_4_58), .D5(mdout1_5_58), .D6(mdout1_6_58), 
        .D7(mdout1_7_58), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[58]));

    MUX81 mux_39 (.D0(mdout1_0_59), .D1(mdout1_1_59), .D2(mdout1_2_59), 
        .D3(mdout1_3_59), .D4(mdout1_4_59), .D5(mdout1_5_59), .D6(mdout1_6_59), 
        .D7(mdout1_7_59), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[59]));

    MUX81 mux_38 (.D0(mdout1_0_60), .D1(mdout1_1_60), .D2(mdout1_2_60), 
        .D3(mdout1_3_60), .D4(mdout1_4_60), .D5(mdout1_5_60), .D6(mdout1_6_60), 
        .D7(mdout1_7_60), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[60]));

    MUX81 mux_37 (.D0(mdout1_0_61), .D1(mdout1_1_61), .D2(mdout1_2_61), 
        .D3(mdout1_3_61), .D4(mdout1_4_61), .D5(mdout1_5_61), .D6(mdout1_6_61), 
        .D7(mdout1_7_61), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[61]));

    MUX81 mux_36 (.D0(mdout1_0_62), .D1(mdout1_1_62), .D2(mdout1_2_62), 
        .D3(mdout1_3_62), .D4(mdout1_4_62), .D5(mdout1_5_62), .D6(mdout1_6_62), 
        .D7(mdout1_7_62), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[62]));

    MUX81 mux_35 (.D0(mdout1_0_63), .D1(mdout1_1_63), .D2(mdout1_2_63), 
        .D3(mdout1_3_63), .D4(mdout1_4_63), .D5(mdout1_5_63), .D6(mdout1_6_63), 
        .D7(mdout1_7_63), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[63]));

    MUX81 mux_34 (.D0(mdout1_0_64), .D1(mdout1_1_64), .D2(mdout1_2_64), 
        .D3(mdout1_3_64), .D4(mdout1_4_64), .D5(mdout1_5_64), .D6(mdout1_6_64), 
        .D7(mdout1_7_64), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[64]));

    MUX81 mux_33 (.D0(mdout1_0_65), .D1(mdout1_1_65), .D2(mdout1_2_65), 
        .D3(mdout1_3_65), .D4(mdout1_4_65), .D5(mdout1_5_65), .D6(mdout1_6_65), 
        .D7(mdout1_7_65), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[65]));

    MUX81 mux_32 (.D0(mdout1_0_66), .D1(mdout1_1_66), .D2(mdout1_2_66), 
        .D3(mdout1_3_66), .D4(mdout1_4_66), .D5(mdout1_5_66), .D6(mdout1_6_66), 
        .D7(mdout1_7_66), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[66]));

    MUX81 mux_31 (.D0(mdout1_0_67), .D1(mdout1_1_67), .D2(mdout1_2_67), 
        .D3(mdout1_3_67), .D4(mdout1_4_67), .D5(mdout1_5_67), .D6(mdout1_6_67), 
        .D7(mdout1_7_67), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[67]));

    MUX81 mux_30 (.D0(mdout1_0_68), .D1(mdout1_1_68), .D2(mdout1_2_68), 
        .D3(mdout1_3_68), .D4(mdout1_4_68), .D5(mdout1_5_68), .D6(mdout1_6_68), 
        .D7(mdout1_7_68), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[68]));

    MUX81 mux_29 (.D0(mdout1_0_69), .D1(mdout1_1_69), .D2(mdout1_2_69), 
        .D3(mdout1_3_69), .D4(mdout1_4_69), .D5(mdout1_5_69), .D6(mdout1_6_69), 
        .D7(mdout1_7_69), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[69]));

    MUX81 mux_28 (.D0(mdout1_0_70), .D1(mdout1_1_70), .D2(mdout1_2_70), 
        .D3(mdout1_3_70), .D4(mdout1_4_70), .D5(mdout1_5_70), .D6(mdout1_6_70), 
        .D7(mdout1_7_70), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[70]));

    MUX81 mux_27 (.D0(mdout1_0_71), .D1(mdout1_1_71), .D2(mdout1_2_71), 
        .D3(mdout1_3_71), .D4(mdout1_4_71), .D5(mdout1_5_71), .D6(mdout1_6_71), 
        .D7(mdout1_7_71), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[71]));

    MUX81 mux_26 (.D0(mdout1_0_72), .D1(mdout1_1_72), .D2(mdout1_2_72), 
        .D3(mdout1_3_72), .D4(mdout1_4_72), .D5(mdout1_5_72), .D6(mdout1_6_72), 
        .D7(mdout1_7_72), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[72]));

    MUX81 mux_25 (.D0(mdout1_0_73), .D1(mdout1_1_73), .D2(mdout1_2_73), 
        .D3(mdout1_3_73), .D4(mdout1_4_73), .D5(mdout1_5_73), .D6(mdout1_6_73), 
        .D7(mdout1_7_73), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[73]));

    MUX81 mux_24 (.D0(mdout1_0_74), .D1(mdout1_1_74), .D2(mdout1_2_74), 
        .D3(mdout1_3_74), .D4(mdout1_4_74), .D5(mdout1_5_74), .D6(mdout1_6_74), 
        .D7(mdout1_7_74), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[74]));

    MUX81 mux_23 (.D0(mdout1_0_75), .D1(mdout1_1_75), .D2(mdout1_2_75), 
        .D3(mdout1_3_75), .D4(mdout1_4_75), .D5(mdout1_5_75), .D6(mdout1_6_75), 
        .D7(mdout1_7_75), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[75]));

    MUX81 mux_22 (.D0(mdout1_0_76), .D1(mdout1_1_76), .D2(mdout1_2_76), 
        .D3(mdout1_3_76), .D4(mdout1_4_76), .D5(mdout1_5_76), .D6(mdout1_6_76), 
        .D7(mdout1_7_76), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[76]));

    MUX81 mux_21 (.D0(mdout1_0_77), .D1(mdout1_1_77), .D2(mdout1_2_77), 
        .D3(mdout1_3_77), .D4(mdout1_4_77), .D5(mdout1_5_77), .D6(mdout1_6_77), 
        .D7(mdout1_7_77), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[77]));

    MUX81 mux_20 (.D0(mdout1_0_78), .D1(mdout1_1_78), .D2(mdout1_2_78), 
        .D3(mdout1_3_78), .D4(mdout1_4_78), .D5(mdout1_5_78), .D6(mdout1_6_78), 
        .D7(mdout1_7_78), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[78]));

    MUX81 mux_19 (.D0(mdout1_0_79), .D1(mdout1_1_79), .D2(mdout1_2_79), 
        .D3(mdout1_3_79), .D4(mdout1_4_79), .D5(mdout1_5_79), .D6(mdout1_6_79), 
        .D7(mdout1_7_79), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[79]));

    MUX81 mux_18 (.D0(mdout1_0_80), .D1(mdout1_1_80), .D2(mdout1_2_80), 
        .D3(mdout1_3_80), .D4(mdout1_4_80), .D5(mdout1_5_80), .D6(mdout1_6_80), 
        .D7(mdout1_7_80), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[80]));

    MUX81 mux_17 (.D0(mdout1_0_81), .D1(mdout1_1_81), .D2(mdout1_2_81), 
        .D3(mdout1_3_81), .D4(mdout1_4_81), .D5(mdout1_5_81), .D6(mdout1_6_81), 
        .D7(mdout1_7_81), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[81]));

    MUX81 mux_16 (.D0(mdout1_0_82), .D1(mdout1_1_82), .D2(mdout1_2_82), 
        .D3(mdout1_3_82), .D4(mdout1_4_82), .D5(mdout1_5_82), .D6(mdout1_6_82), 
        .D7(mdout1_7_82), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[82]));

    MUX81 mux_15 (.D0(mdout1_0_83), .D1(mdout1_1_83), .D2(mdout1_2_83), 
        .D3(mdout1_3_83), .D4(mdout1_4_83), .D5(mdout1_5_83), .D6(mdout1_6_83), 
        .D7(mdout1_7_83), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[83]));

    MUX81 mux_14 (.D0(mdout1_0_84), .D1(mdout1_1_84), .D2(mdout1_2_84), 
        .D3(mdout1_3_84), .D4(mdout1_4_84), .D5(mdout1_5_84), .D6(mdout1_6_84), 
        .D7(mdout1_7_84), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[84]));

    MUX81 mux_13 (.D0(mdout1_0_85), .D1(mdout1_1_85), .D2(mdout1_2_85), 
        .D3(mdout1_3_85), .D4(mdout1_4_85), .D5(mdout1_5_85), .D6(mdout1_6_85), 
        .D7(mdout1_7_85), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[85]));

    MUX81 mux_12 (.D0(mdout1_0_86), .D1(mdout1_1_86), .D2(mdout1_2_86), 
        .D3(mdout1_3_86), .D4(mdout1_4_86), .D5(mdout1_5_86), .D6(mdout1_6_86), 
        .D7(mdout1_7_86), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[86]));

    MUX81 mux_11 (.D0(mdout1_0_87), .D1(mdout1_1_87), .D2(mdout1_2_87), 
        .D3(mdout1_3_87), .D4(mdout1_4_87), .D5(mdout1_5_87), .D6(mdout1_6_87), 
        .D7(mdout1_7_87), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[87]));

    MUX81 mux_10 (.D0(mdout1_0_88), .D1(mdout1_1_88), .D2(mdout1_2_88), 
        .D3(mdout1_3_88), .D4(mdout1_4_88), .D5(mdout1_5_88), .D6(mdout1_6_88), 
        .D7(mdout1_7_88), .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), 
        .Z(Q[88]));

    MUX81 mux_9 (.D0(mdout1_0_89), .D1(mdout1_1_89), .D2(mdout1_2_89), .D3(mdout1_3_89), 
        .D4(mdout1_4_89), .D5(mdout1_5_89), .D6(mdout1_6_89), .D7(mdout1_7_89), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[89]));

    MUX81 mux_8 (.D0(mdout1_0_90), .D1(mdout1_1_90), .D2(mdout1_2_90), .D3(mdout1_3_90), 
        .D4(mdout1_4_90), .D5(mdout1_5_90), .D6(mdout1_6_90), .D7(mdout1_7_90), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[90]));

    MUX81 mux_7 (.D0(mdout1_0_91), .D1(mdout1_1_91), .D2(mdout1_2_91), .D3(mdout1_3_91), 
        .D4(mdout1_4_91), .D5(mdout1_5_91), .D6(mdout1_6_91), .D7(mdout1_7_91), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[91]));

    MUX81 mux_6 (.D0(mdout1_0_92), .D1(mdout1_1_92), .D2(mdout1_2_92), .D3(mdout1_3_92), 
        .D4(mdout1_4_92), .D5(mdout1_5_92), .D6(mdout1_6_92), .D7(mdout1_7_92), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[92]));

    MUX81 mux_5 (.D0(mdout1_0_93), .D1(mdout1_1_93), .D2(mdout1_2_93), .D3(mdout1_3_93), 
        .D4(mdout1_4_93), .D5(mdout1_5_93), .D6(mdout1_6_93), .D7(mdout1_7_93), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[93]));

    MUX81 mux_4 (.D0(mdout1_0_94), .D1(mdout1_1_94), .D2(mdout1_2_94), .D3(mdout1_3_94), 
        .D4(mdout1_4_94), .D5(mdout1_5_94), .D6(mdout1_6_94), .D7(mdout1_7_94), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[94]));

    MUX81 mux_3 (.D0(mdout1_0_95), .D1(mdout1_1_95), .D2(mdout1_2_95), .D3(mdout1_3_95), 
        .D4(mdout1_4_95), .D5(mdout1_5_95), .D6(mdout1_6_95), .D7(mdout1_7_95), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[95]));

    MUX81 mux_2 (.D0(mdout1_0_96), .D1(mdout1_1_96), .D2(mdout1_2_96), .D3(mdout1_3_96), 
        .D4(mdout1_4_96), .D5(mdout1_5_96), .D6(mdout1_6_96), .D7(mdout1_7_96), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[96]));

    MUX81 mux_1 (.D0(mdout1_0_97), .D1(mdout1_1_97), .D2(mdout1_2_97), .D3(mdout1_3_97), 
        .D4(mdout1_4_97), .D5(mdout1_5_97), .D6(mdout1_6_97), .D7(mdout1_7_97), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[97]));

    MUX81 mux_0 (.D0(mdout1_0_98), .D1(mdout1_1_98), .D2(mdout1_2_98), .D3(mdout1_3_98), 
        .D4(mdout1_4_98), .D5(mdout1_5_98), .D6(mdout1_6_98), .D7(mdout1_7_98), 
        .SD1(raddr11_ff2), .SD2(raddr12_ff2), .SD3(raddr13_ff2), .Z(Q[98]));



    // exemplar begin
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_0_87 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_1_86 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_2_85 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_3_84 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_4_83 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_5_82 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_6_81 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_7_80 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_8_79 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_9_78 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_0_10_77 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_0_76 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_1_75 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_2_74 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_3_73 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_4_72 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_5_71 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_6_70 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_7_69 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_8_68 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_9_67 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_1_10_66 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_0_65 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_1_64 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_2_63 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_3_62 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_4_61 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_5_60 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_6_59 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_7_58 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_8_57 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_9_56 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_2_10_55 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_0_54 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_1_53 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_2_52 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_3_51 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_4_50 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_5_49 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_6_48 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_7_47 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_8_46 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_9_45 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_3_10_44 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_0_43 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_1_42 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_2_41 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_3_40 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_4_39 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_5_38 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_6_37 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_7_36 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_8_35 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_9_34 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_4_10_33 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_0_32 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_1_31 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_2_30 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_3_29 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_4_28 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_5_27 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_6_26 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_7_25 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_8_24 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_9_23 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_5_10_22 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_0_21 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_1_20 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_2_19 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_3_18 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_4_17 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_5_16 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_6_15 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_7_14 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_8_13 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_9_12 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_6_10_11 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_0_10 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_1_9 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_2_8 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_3_7 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_4_6 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_5_5 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_6_4 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_7_3 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_8_2 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_9_1 RESETMODE SYNC
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0 MEM_LPC_FILE pmi_ram_dpEbnonesadr991416384991416384122adcc5__PMIP__16384__99__99B
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr991416384991416384122adcc5_7_10_0 RESETMODE SYNC
    // exemplar attribute FF_5 GSR ENABLED
    // exemplar attribute FF_4 GSR ENABLED
    // exemplar attribute FF_3 GSR ENABLED
    // exemplar attribute FF_2 GSR ENABLED
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar end

endmodule
